--
--Written by GowinSynthesis
--Tool Version "V1.9.10 (64-bit)"
--Mon Aug 18 15:51:03 2025

--Source file index table:
--file0 "\C:/Gowin/Gowin_V1.9.10_x64/IDE/ipcore/INT_MULT/data/integer_multiplier.v"
--file1 "\C:/Gowin/Gowin_V1.9.10_x64/IDE/ipcore/INT_MULT/data/integer_multiplier_wrap.v"
`protect begin_protected
`protect version="2.3"
`protect author="default"
`protect author_info="default"
`protect encrypt_agent="GOWIN"
`protect encrypt_agent_info="GOWIN Encrypt Version 2.3"

`protect encoding=(enctype="base64", line_length=76, bytes=256)
`protect key_keyowner="GOWIN",key_keyname="GWK2023-09",key_method="rsa"
`protect key_block
jK05pR8SRRPfLSWSMbIhLl+a/VOzEimTQh/0YSOlY3MUVz7bA0rmwivVU+To1yzMDELuH8Imvl5w
gQqTTBbiFpnKLOyYA9rHDnETySSG63Vn5ehfULZY2AqUKMZUdDNtwqDKQMW9vfS2wbJ0QNMW/kJX
N8QrPKAm6KJzZ0btzNfFo1a5KInm7v50RGvICvqJWSZgZNyf4AeQ+vU8UqRS8esyhaSqNxZAvuQ9
qKUd9jHUlF7BjNYxkFcutjj6Ms3jAXwk2s88iy6bgI1fACHcQN4MCYxRPuzRApToDu38epcOGcr+
w060jyp0hZqX8ryD6FqMj3Ubo5U2AB26o6HLmw==

`protect encoding=(enctype="base64", line_length=76, bytes=240224)
`protect data_keyowner="default-ip-vendor"
`protect data_keyname="default-ip-key"
`protect data_method="aes128-cfb"
`protect data_block
3YFOrHLypeJczoQz4hF/LwhuZk8AnQ5Til/uc3DjJoyVwh8RotSycU62iVq8jUchFwmGu7fjHdTE
x3XnhjIQn8xSsFb0dooR1qoxq95f3oCmwZ6viypsr7OP5r61Z02GwMdHGz9/FiNHSdusTLqpswNM
emeEaV1hKafk2al8oAppAvZOY1JEEflQn1hjA0FJyzf7O/KsY3Ork5eKysbeMfvTnq5fofchXCZD
8WVnsDwOCDGUYcf0zRXiIjfLRZaB/YrDu0iJXeYxU9Zfs7AxXz336ShH1lgq3qEKila6qa8aeNk5
BrvAVPqmyT+qGVj2Nqc+VcF59zrXLKncqJvWRnqgexEk6LKM8yjktxQmmw/6pFZBuNti5Ov3w7VG
5RtgEaBtK9G7QWVlAne10cbFW+vAAPwFGrXmBpMQH1JakZ2QY+NYUxLwlOIoeMHcZ7Fz3k5VsUUW
UbmlslSiVIR9SqXrkufcoWpfxHuMkYWQiPHIixRsp+Wo/MBMP+hF5Ci3yFrQdc5ZmS31kvKgLLNG
zx8a2BdmwEgpyOZwxkZBEOyOIaDNd3AVzMdTctApFGsYSAXaL+iqrZ/DpuoKLCwyi24+1QvnrxF1
4PRC6x+oTwRKgN7wf2vBk5X0kVi7n7qqLyUYmFirF0kafOAEF5BirqlY9NC7x/k3+F3/3p54zg4D
d/5fkRdOuRVQRapKnuel5cgjEdADvK0m036Zpr9WMtLY0eAiDavI1naWuuC8mWp22M9uHCDxAXfH
f8ZxvLWexhNWcX+CXFXlwOAMOY7Yr1PxSOvyEmvupZnl1z+Q4EB9oQBp3zfQpARoBX3NOv6Rl/zC
WV9KOfeAs9DywFPBBGQrjnfalHnKcQrMhta7H9xj4cGYJvuVQWfOmSU+6dtLShLI4nCg99vxphmk
d60FyuUMrImggrUZeCLFbyRbzxYkWy911y9ZOEslRGM7mDolgw3pCDkXAO00PAyl1btFB3eBUMJL
LCthZexiaMvrFQ0X8IE4IC2SVBQkSm72Ym0U1QNJEYmoGxlkyd/R7oISPqXiVBpnv2hd4fsLY7vj
zwFnY0SeU9CDAT+vw3LTNkNxZkQXrZ3CWKqSAddZMY0+hOk9GJXjzWxdFkwaV2fVbTcMNn1mClNo
3Xu/pTPXZJCij3ESLkDr1u7zaCjqSRExGc1EUMB86FwvYUP/0t591EmxLWfl9uMifkqjuQcSje5V
bL8zu5STg9YOdn0kpndLQdd5m2J6yynI9XMZHeDcBCDwHby+JnsCggRpw7MgFvjncUkoykKKAPcV
wrctj6uEsBLiH7ZDxBZB4+mwNdThhthNdwpgWG3D5c1c78+ktRZ7yZKwa7faxonPasKW//CK4gNu
mHYzcuonHPPmiBpF/VfdTP9P4AA2/IQY6yCkcEK8DThoXesZeM+IXEF6me/yesIiM1kSmjQNXKBh
bjzruIAlRSPeeLPG6gqzRo4fJZb61K23xYsnDC7Sa1Q7HJMqwgk6NLNHWZF5m1EZ+bmnrtw5rch5
15QHNVm72iHA4gfVpzxXRuiQAhEGWYFBMAU8oKao8xuUK29qJqfkAzN48ejZEcD23PgPbq5NsGOj
Z4qrBR8A8zKre0wG1KbAQQAW3o8apJE5PNl/G6pYTbL8tvn4SMRQFAsalIO57Dj3Lmm+mvPIrTUc
Xh41gLJNNX1oVRH1svaT3wMUwODWTgs/71H8CkAztbHxvclS4oDmBHRXxhj3etUG5+g0nowzmul/
UStkuFpQCFhsA4uJaqeWBIayhuSqa36683jdF1BL+mqA5IYNJTH7fZLk/UmP4O1bJIrn7qpzJubv
b+cH34u1z4FrOdR1xWCk6z+d/FaOiv+8rdeHY8YlI2hwK2yIW7Hu3j/iPnZBHAsXvPrRdsEoVXj5
gj8T06JeASSo+hjB/JOp3i4H95OsgRVrifdIQhqUMRlflpD7fbZPcPvdk+BmTmJ4D+8lNRpYtnwP
2LcFMectrQeLO02w/coUHQKLAvwk+29/pMlPOrK2VB/7mAXYYPwPSghMW3NqjGa2UlrevhctjKGp
tNZnDJNkREVY0hyNrfrBHAM4gVW+AJ+Hu5b6XsYL7gKmSrOvD1lnG3v7JsVxBYnx8StbnTYv5N1+
JaAuFKTA+mvCOO4Sc27QY4MXGI2Dix05u1YTDwvRT0mS2y/+dhyKdazkGr2e3LVhowW2+6h2uG7H
fXBrB7GiV8bYHbeWGotOKpuGD/BZKvphanreh4xbVndEZUjuQ2GUBUdp9Cmcv6bVsFYP6GWfz/Nq
/1OvQyfvPeu0N5Y2Kqi5CNTXjtYzOdmVWneUJpvKkGYCtMYVl/UNmc7WBjBmXK/DE7Ipfn8Rnd9g
K+0umGhMUyeMf6K+7tiF/t80i1E7AhcEOqAyzOop1qJNJWJDzq/DBRlBXMH6V6ZfwbhNXhFWgDCd
bzMwyuxFzbAuEtdXPA44M/xSkTbEf+1Dml39TIlBuUHKcrpQpZIGSxp1C3Pqd+00y8KVSa+GGZpS
zjwzq1GP+KEz7DzpnnaL2JKDrYv8BhoKV9nhC9tAQg0rTx1clBzB4nEJ2EilMJCFJN/U1pq0/71l
RlQbpfnCMW0hRnirA+vuDLR0hHTWXkgbGXJCSvMv+l+5Mfo55TB+37Sc/CMucCcavoAS7fEC7G4e
6xRlDePVuv12slICNKA+3wQ7FVAfQdJM0oi6+tD5JwxmOYFCKjBjeCvKCANf1rHWTLrtLhFtuoiG
dXQarWMuYagqqBn0TlGHVWiW6O6Ynmc2gzjyCwuIqe+qKUwNiuAF8iF6DDLzvA+vwReRQyjfBwsd
b5TZBKSE3GAS/XGaxAAk6XM2ABV0XHnR05jAPS6ECjTNhFvupHe/scp9MchaKsMlvc45yP6l5kLs
5JFfVfOXv4AiINkS6t9X6PVrHlFry9S4cr4V36H2sZQelW2oTtpTbek+nfgu1c7Ii2O5Ulf8TZV3
PscZ92pHPL1cwhhu4QmfFu8WOZTNueUuVTkNg6zU4rBwCj62lNJgLL/jiG372huRybBcu1oKsXoY
C3VCBJ6nffi9INenSibNCN5isGa6HsLExabAr0TmS5qnCQFrIYNgBAevTdnFtPBOW/n6r654RhK0
ucamDu52kJvNc2GnwI3Bnx/dCarZs3Nu6DIif3bBDceo4DiNlg6nHcE/642xKrQScZvBeEdF2tjs
XUDLf8IfMyryif9+W6zwBiJzZtC699RwbnXz0af28CJpg8WbnDL8I+uMw88xKhjFAfNGPVDqgpdq
1qsxl/iSAo6nfE26wXtnlo66lS6zLakLIM9RYI0zy2oaPTps5LfQYQuz9H6YYPZxg9DuGM7Hg6fL
Reu+qn7tdpdhjQ8SdPEn1kgFxz7ns0FkwisHmwEYlWrWmwZWJbKpHu/dfRlsSh1hwkqzycXFJISr
6Xh9ynlJCus6w6a+O2U806oHcLyXtDfVpNnEil7hlkxQ2iFPqoRazXt/rAux2QFPXkWBfFKPJ0om
UYYIs1Iee7xgKjofrXDYYxL6HjIKu6NR8JH88psABnQx7t7OEkvlKYbnjGuPskC1UodGau1B9Zrx
r+MJ6ST06syDBh0vK+7RHaUk3mDXD1sHn0UB9peQBCxv8gmFOzvlg4AcdRDWLqkHePT6BlQgghgq
H2XBpT0HgEhBJrNB09blJiJzzXi2QQiqOAoc1CkWTpp8Y2AGOXEXOUS6kjJeTBceGXjD94pmyX0I
DcqtR8AZlhnFcmtU9lrZsKd5KMUZqKhCdoZ5nilWrW1Zv6jbK19LGtmm2M8lgMPHmonkEbR3lB2j
2c+SM2pq4FeghXi9eeMP8Mi6T/7zWXSBbAlsjrhYxU7z0Vl2UDMuyPVXskaJ7dErG0FP8NmsuVSK
m2hVgy+u58KBws+9D3dQ6AXp9GBKFYp3ycX9D22Nd8XT7CpsA2hgi6fJhRRDrEic5NYntpB2BjGQ
LkjR0Up6IzpociQ3FfKotyUwKWIQYoPA5/fDWvh19osdTpg0TBdfL2Gx0XNX/nm4d1ZPg0JRIXMd
2cJ9Jjo3V2at18xYde0ETK+P4xRC15kM8tB0q3enxWzCKxnWbqxlVJasTl1vq4+KGu5OwBp5J4A1
l4YzwiQpdMDfjaGaMMMuMZLd1hghv4c6yh5suWyzDB3Jra5mLwE6laHJG9fYXxTp7skgvxFPu4jB
QICsh0ayFbgE1XMNuKdrbZ9QrVI39fpmi6aKnJBXQW39AaBVbUSC5psx4XvlfmiNSHPFKkC5VQaU
8tysXwzrmMMF0IpW74qVx/h8mLu7PDX3s5zCJaxlXopXrCUb5P9SaqcPl5apj946or2EVJXu4rf2
jZdGAvTmlAu7W6oe/kDWMLFsc/n0Xhco0WKyYZIUzK7Ac7pTyxdiKWMON9XpEYajw4VftNrKs9YS
6ZPaiw1O+chHDx2lbEnbn4IsdfL6YCnARqu99nx2HXIn+m+/7jz5E2yaQeymAw3xzG7JZsQ/7s21
s04rJ2o+j4ePK5qUy132DBbc6jNecc1+EhcoecU/ObsMpK72r9ulfrdB4EPcXHiwcnovFRtJSl/9
YLzmD5lVOaQdz9slz38vC7gfFWuP5FJMFW+RWLQc64OLG4W6ni5LrqLdRzZiJE9x/DDw33B8FfsP
W0t+UJuS0X2E/h3LQRQdIoDadGkDH7PQcQuZCkcLydXFJKZMN40nLDMXQJSx3/KfSyTBLtWPJMau
xlft5Xgb8ehRmAkvZ+wbmfjtym2R4DRRGG2hNTWn0ohrS965XkX4kkKNWaTqLXFcF9wlI1nSpfkj
2KplFDerybjTBST/l7QJUZHF3l7xkVqmWbtG5vabYVe20aPDIB0DIOOBgSLC5rW472bxmeZEphtv
cd2cNsx+R++8vlTRII4Xo9Yq+2q3+R5QVOZSx3f0v/vn/Y5/m8/yNhCw5LTXtZEtO90TzMDSUL6h
h9fRStpfeRfJ9gD4yXKmwACAENGv6GktkWTY3Afoyrb9Fo/CL2fLNYSBsmuoEUFrJ0fBhL3Y1Vb4
VSEpkrhOB4CRM9gxf3yesNtRfFkpTdYMH6fVAAzkwtRS6+/5YzdoJ3x1QuChv+TpJT5IM+aL6JB2
VcvhBDpIkG24lLaTznKiCdd7IfQDjd3l9mn/y55gbdpSg1yztqMVjHqwfYhiJezgVMaVS4WMwj5E
PzCSUwvt2ppHkD2e9kEf30kjZF0BKocYTkS5mNj0m2FAuhfplbR9/9ta3KqsF14j3VWGyDgpcQpz
Q7ybKLSjoJMY/cKjw+Q1VYifv/oVHM/rfbOSqszpphUGhRQGnp/74S/88SFTn51w5gOVKC/nB3W1
vZa6bNFJTL5Wf+55oNsZ7L65+4hLc9e8cR4OZ+1Tz/ftBgNxXbb9CsKkgqxqwICLwfCc9GN6bjrp
a5i/sHkB5x+mnuB8Cv6mh+QwDuLMf7DecxT3Yc3S+BdHPkQ4zSsb5/dCGtrFJbHx5oCBmNichwCX
srwF2VBcqKX01EYSYryVrqKHmR/sTvTQ//pdwRS+ul6tuOxcBUB1M3I+tgAd1kVFWkA4XlKO9vMc
bpSVBsNBjjzZZHzYzfvOO0nkyvwSrXQuMrbhKlcdSbPHVFw87piSENcATUEo4TqepaLAxLDu0tCj
vLUGc0U2Wam/MtdHyR/Rp2Q6eyL6Kyocvle1H4oA/ENdoUpNuKWawrQ4d9+Ls44uWprNYx9OPEIO
3Ju5azmW1earixjbWToyT9GY1T4yN80dF2pzaVkypAfsI3do1X6+icF4ETpTUpcBEHceaVU80cjM
3OpFcTjqCSsR3/8epU20AOVP4hI3lpqu/ut6eSn8ZtPm4T1rr69Ss3DIjfy9qOylHI01QGOriR6Y
VawfoDX+odGlAXOK2WLXQVaGV5r8SazHXvpCixYbBVTsgoaoQsT0ezK6FtlOewN4GJm0xb5h1LJR
cgYk/mInGBLbeCflYvqylGCjD9mGe6gT88fBBn6sx1/pQVcb6wn5MUss1WvMwkMvMgA1j7JQWNFT
igrST6UxSgDsM1SFms1k7u2aXVIMPVX1FNEsJZ1El5Ghi3o4WrTEMskEZ1rMoL8DE5UPMd5cMr66
itUxLq8dDDBwprdXTITzhvOfh9rZ8TppBLdywGC3AseYIS8OU3/Y8ZnK0F42FmRny/cUjqsSYwoR
hPh0ua0q7lSuwLLGR/aqNRWZssWw/UhmwnvQcZiFl0HR+oUoMcWTtOyIwPMKWM7Q63v1cLhHroBY
l3XUAaWvlFIuah4X0Sas9I1LACbPNsm9TnGNBa7Y/gJL0ME73lZOHEmGjrHX2eyCvqXj0ltkqslJ
ppT/U/CBeUqQDqCosP4QJspaGKrs7Zciz4rADg73BOcqJDpnd8SThqKsXGhCH4tuYg2AqZCjfh5U
bCLe5ByGvykGAAydWek5R1D7Ysxl2nMjCoLN1+HyFBTuGM5FjpodvaOaWtDXn692LD/20jhYbPfO
EPtT0gifwxpjHbo+z2WucFu3yunXJO0SgegovmeowcUSJWAzkmIzk2uKhwouomjAA6MI4pKfD0F4
7dtJM/a2CxNPBv1KTbAGKbsD3n8MHq3GAhA7XNMc3BoxGbNZpi9QQHIk+suUfTs42XZnhonveCXt
dIpraKaq67xBob3uL1+aX3zzo5UzcZisriMKe+llYTLbtwh6Cqmt0wvSiu2S3CPEYYfOPH5L1grl
9FJoyVRQsifyUNX3/Idh0BdtUCz9tvuu5V2iM6GzP2TuKq5aySg1r+v3DA0pr0Zb/Z79DulgZ2QG
mg8rrl1Zmh/Otf4sjf7E3fhql+ojpMjpqIP8bhD/IhyEkt9fzNeY/Qhs9jXl9GBVV7PeEtujx6JF
1TJCWi/aK6BUFQ5nYs99OJS/d1mydmdKuuLw84pScsbaOL7VIkKg1HCUzwIv3yRQACRAPVNN/KrL
IQ2iNymqcMrR1Uzf7HVFbmVlqdnzrUc6W8v10Y4ajEQPQFQQl3if/8twLYhwC9suiPzghypT4O3L
gOOhmYKX6DIPrmZbmhtFGLOHw2mgmt/hijpgcX1QR7gtW9o42KDRKbp/hQUgwhEmLuwm8pdmAxfp
9h423OGvJ2ziXo2YPSgBYHtzN3KIwYWE2E5c2Dkk1gG0DpH9vAr8Q7/2d/Og8oYBbkMnemvQPk2K
n70HLYCTf7yToBVl09gOu/cr7KCrtdiLRvLImXhNzVG1H06MQ91HYNHg6SN1b34W2ofgEytHc3l6
jFm0z5/nTLR5uyzj8lIZQ2R9zlN5/TX7K92dguHyLxrG25nZmHwUjxhi4xmPR7Wc4JmbLCygwDJO
RzhBgpXGhEy2LrxJzbcu/syaR/8wE3yjLs5K3kNpsRkww5GR3RK3YxsCfMGnjgCHkgl2TIPCJ4ab
NNipumbmtWpx4c7JuXONQDrJQMEoVHfLKR8v3ECIl7JPcSuxYIXbpvtPXF9seYP4k7MhEYOTWr8Q
Yr4UDvD4J4TtE3SYepYnTNrk8MjXi8eLz8kJ9c+EBOgRpxWhdyMLbE+XxLro+ewYIombDWlH2i+b
J4BP20L6et29OpO8LtSnm8XUe+xZzM6WdwH8Gb28+ZPVpX8Sy75zlxbZvYM4I+7FjyEgO2n7td6L
aQpzDG0D1mkO7WflhSBJ0zV7byAUwYhFdpklNfw7ahmU97yoAQl4hhw7U2SQ3VmST1/w4B448jhS
4F5muFDvmHl5O63xs5G790JB9m1Kd36r3/C15xxQznGz2T4r9RovxU8Mc+RmiCsieWCLX9jtR/kq
5+lP7sYmw57OzIt3Fu4vp9dhbXEh+LZxKNwwHtxu/TqeMGHr05AgjUxV7tXbN+m1W+L4XKGfHAYp
GeERX+85vqCfgOvn3/iYj3qZl8r+5N/W7DrhC/gQsyzaXmOH5rwFBqMsrPhF2Vy0Iebjp8QQv01q
HZ4F5ZFyyQTgP2HOptN+oVWPyD20Y2f0nmkISGbuJL10iXrXB+yJm6cdY5HIQa8JOds9e7TGGy10
qL2JM1F5aNqXiiRxYQb8+437D7ehEWv4qsDtzQS+cDiVN5Fn/j4Ar6IgrnMLU8cqgnYS3XBmLvQE
KLg9CxX/hShgB2gYk+nIiIc5o0F0eUpJr5xxFgpO09Zq1kBTCH2UQdIqahzbLKHHD51gDnDKYqU0
LY2bO6NuveHplnDpBf9HeSQ2acAbXnD6l144J2yIrP6Wy3cwT0KGEnjFjkWEhd+mvt6bw4jy2Z4N
VllHtJ4CO/WgeJ55PO22QPXr7ag+5gmtjAnwEOVJdKQwz2KmfiLDo2gVq6U18fukW4Ym3QCmoi7j
ZxrFpMumSPfIvLwMqBy4/forsD2i+TREGEZVXw6+U6CwTCWB3YPSilfs0YL6sBdwhAxJ+ZjuN779
TUPJHxIYv98MMbNHmINtLWRj6DbIBcHxW+/8fIROjRRsRKbuKGXE5GI/hBehtTn8FQnGPGJ6fN56
h0YTZGF1Nn7Kc0ETfbjmuaUxPOXa3YhnY/qmVRwGBNYXmBOItlFmqI8jVKXKDnYeEz7NVvMh45sh
aBJf4zAkCyJSoIoCyvomPLOkMKvmTpWnQ21BGgtii/Guo9+XkWAMxqBXhoyWZ46yGzLjamdOnvIL
0kEbcZJaoDCT/bEUz7hbxgBsDJjYosdJfVUZOKfi0qKURGQaSWFxg50Uuc3aabn6NK8sJKMnCu84
R+S+OlSwsRKoaT9yM/fwfD1Z3ewtLWWJyg7a7xnoK+ewKVB8+UmgfMHs4yD2yDjNvNhD9BjqK34L
DDJiPB97rDSa73LZbsilcQhZlHQ6jI22Lg7tqlqXMiXvnKj4Jiy4e9OqpsqIbqA+xLIXD19b5L1c
pqFGWM7M5iJpAi1klplqEU1/tGMmq6yaEqXTl2X0geR/c6Qyez2ZkVnyyVouWTxZzr70qcpKZjzn
RO3Lf1lx+T10t9AUGPl6Ft7cal9di+qyig1ZS4EmDPUj38oSRNYq1kNPbO9eD5xZoootb0Bc1F2j
nqm/zYrp6gLiEcRC7aUqjKvovOZEALuRDHPOJObd3kXZX3otnbsmT6zAdkh/M3szfh/nLqZzokkV
SQU/aeYou+g+qHFL1Y3bDW19Rih8sWHUX/w5sVJvO1YjTf7vr+KI2sNnEWWuzb6z7nrDb9IlNJme
ZoF6Kl/kPyQ5IR3PxsY6VWb0foOuBFovO8MRO99HmZNKmfewi+nB9K2gsiigQK3VDMq0Pb1jLMWf
2EsDW7weMBh8z8clAIiy/dTYsk+OU3SNC1WCz1qPulgESrieI64EVyEKa9qyTB+/VD/EIT/EL3Lf
xxZNbYcmoVv/wELuRuwo3yaDh+FPXDXWaa3DkrakWAJE5dxYN0jdpJsLdDEz/noCDGRPRTwsdzzu
hbfS6jrzfbeCBCMOe3ANbchImsHNOIJo/xDW17vnFtwvm84dmhYaYNhvxTnXY69Y+0btYKUPxM5T
h8dtHwduLe9wq+0bgLdnctw3ojc3coCCUEMAsxjQShKibE8JrJG/jshuHW2S7GGs7A5haY9ZcHs/
7jzmYXzoXIO0qbmW7U8cYnnhuzZYeFT0aMlp7t9cA6WOnlMg83biUnkGvOCc7x/4FUFyCyNBRpkW
SI20Wn2jl6/gak0oVdceVw7+R6Wtu3zUj6a7CAzLVdoF5QSlEo7FozkxHHU1YiMb0kMW/zLZvICX
JTlEBrTNC4s854tzv7eXLKCyCGxajmwlq3l7ukd2yLTUsUvzFu1qlrgcxD5R98yLEvNE7LGIENr9
bZeZNUTIGXfV/bOHzQHIZR2OJvbMiU785nGb3W7biKRJhwCjeQksj7XdB5iTb8gIjez617PR7AzD
yyjusksOCUL8WDtgHOCYVS1CLUILRb3sRNTK8jTNCrMRaEtFFioQ/DnLXzzJ+NyIm1TmVkGWLlSh
b3dUnOb6vWBmUhXb1w3xXomVGi71Kj451CG9Q0ogOD9Cu9ku2XRZ71Nmu0UTECPNU+ggtPcWBEqx
yfDYKtF96fUd7YVmH1cmtc0kfPRMgJAQPHdW43Urp2sH7boNEOPzg4vzVMNrt+1jLlRCIwUozvTG
RuPW9TNEQhX4y4dXufFoWx3jOlMBOJlVU3P585rT838CA27w7/ZsgUC3T3JcgXR2/0VyCKUtNXS8
9j7vPNMGPAHpa+gITiABL3L4q2/VQYX3DyQ4JZVL3mUYdqbIjbu4b+3KBivgoaWEkqrtRTP+8nui
SuVuqIToHY3NpKBGUuMDOwurBGKn6RC1ap+Pv9zKnTgiSAAzXhJTrTQcY0ZStD92nZR8YfWWpi3I
pVgkIAOauLblyOgDUNGR99Gum1Lif+bGhYjIE6+8R+svna0mszlN88QWoCZg134TymLDr5r5AZQA
XF+e0cYRZA0n1yNaWwedYkXh0Basb9R7SBeIisfhRgwxuZQ8seky9tqp0k6FH6Mh2aDuUaIEgorM
YPSOMtXymwVTWOlsLPWH5D70uYNUZ1c12mKHViHvNib5ahifOTX85daR6FZIwlchxBQXfvgCNoYl
IMoGo+B8irxWdyV0aQ90u3WEB58SaSxKzpKhCkKDKC2ntxbvWSffX6KRkm1CKL9Yzz3bgQtOkINR
3eJxQg6YsMFvqI2ya2fT/IKqoUPdfHCPsqjpml34xlDhuqmY/RqNrElWtR7j6P3TezUg0OyY/HhC
v5hbOuqyFUN/cqHXwzVt5+bBIKq5ynW0VyEIOxNqhgJ70pm5U9do1xWQVaBxfuMWOb60OgLdUDYC
KcQ45FjevOl3K5yYAU0BeRvWD5n8hQ5T7ZUZrl8/QqV7EI7E9otW75P+t1+EsxkdoBwnhMF5RymT
m5g3T9wtW4SjP7wTG1O1wRLzdRhtJhboMQx9yb2stHI5fwBYH6fcp312FqfCfTdVyW2IWAw4VD6G
sB53MJCuBJAQeD7Rd8HZINkS1rd2RIAK9zxURIUVReP1l9kN4fVUdolkuS/72hbDSNHNCOsLGSva
Uqso5mF+N9doHfwFkybgraX+if/sAJdCffG2kkTYAGVI8oHUy1ZMxKpmWLIT3m8OKfVTjbZt4zok
8iegqpfTWFx15tjoJsQXX02U/mnmDmKqKYx1v39Fh+ChsnvIcKCKf4tx9yo2sH5ziS76t3ovaX4q
m+SF0lYWzQPSDW74G43Ilhl1htnIP6KybPWT4k3Uh2VCSWw6n03JNcKvU2oF6ewqGqUmgKBw3Vsg
u9Wrx19LexaZUX2iWD8TrrXXuCp9XY8y2eDj5yR+JMWdCVSOAAIS2PAn/SCBoGuXXASZ3+fEz/sS
FCp/ZdKYBDfuVYIyrrlPWNPhaVS41pYm6ScVE8ghICjoZ6jWn5Hph8mM3Gs/VgJeuDS6PkNTbMq+
AU+BF1vkGfyMY2tzRpWqKuhOIux/tMx/AcGl4ZBggrcf7Ppr9c3lkegX3wrH9yojExwpY0RDWR+L
NxHAUJsZ+eRXH4ATOh6DIqCyrYqZGVvHJTvxym1Pu3pXExwXAJ3Vmh7LBx1moTp10pETuVx049l5
e71ssexulEr6TgBMkeaGVp+M3aYLh1GXfuRQ2o3qXCxG+l7RifZz3pNi2XEmu2vEsoIjgqeTUlEA
1iJKQx5iUSbjEcfXGbHsWbXlq3jTh/9Rqhm8IZFzY0z7KL0RaTk6OBVABd7wkfMcB4AG1DSJVacP
4Bh4WA8cv14fQvKa3xlJc7nObHf1BScvF5of3CXnKJWLcLfSpbhw6xEtXyZQeIgj0dWuc/0fDU/s
43dzdXiFdJcP7byrSpeIJOAmB8bDQ6DEKuRbOUf9FYpe3hrscB7u9rAGo/NTmtXpIssk1QxY2sH+
kEvaJvg5jbA+HBARvorQ/q/wMa2H3Npxjnykf9FTRKsA2psSedp+dgUPGTdtZZtbWHHl6l73TQAt
D7YmD8dP+L7z4ILgPE3ez4qjE03VB7/Q2kd7L4Lk33a4/yg/2R3t7bU3CzzyqR0YMsIZQ9HPtZI0
KgIIURbkyzuTa8oT59w9RIwGEmQChW7u9oTFWRqZd83aLRGRr8TjJWyMtJiALa5+vHMjCPS3+jpZ
Es/WlGD+bObeYtgNXpQ2PaB9FPfL51Ojj3yvSTmiJgdltkeLA1EJ8YSdx4mhXExKwOYvjIseqr5d
1vEcEwCOzyC8hiYn4jbw9/Ufwd6CcUSBcqGijoQtdTXhQwwYXbYlam+5iAY201XiBJg5tkewwvZl
YoM4fMcUEa73cSicvxMMZlS43QvkpSVr7Bzu9+UIc7swEdAkqpZZnFNJtOBP0louVK3IMEzyPAA/
Z3Gm2fMm2hW8bQN5jQi3uDi8K4BPKHxbll4ZUjqe3k6G6M+jk2nQlLphjVQX3C3HyMv1GD93J+nG
EAnFCsfOk0tHa5p6Mq9Zv0Mocp5MGcvoVKUiNZ24Op4cglhlMV5GCc8rsOsk7IBEPgqHD52Cl8Py
vFXsPhuEbbojndXWshqzxKUZorUBam30Hq0DLN71P8geT1hEA85e7jrrLjE3Lnp+gnjW2Y4OgO/l
YktRA27SG//YHQSSSAfhxpx9LGVquA2XT8LHfgAhX6j5qPLWgctqTqCeOP1JMUWqpomv4QNPQphW
O+cqDNAzsP5WzlB+zWWHikO6IWjQ08zjHzk5wNCxdMsl1G/Vy9/6ofN1bQ7eGHt/suXWEktaowRR
JPr7KtFCw2ow3pcQcKf/SYSW1OKuJ4dOz06l8O3ToDgnfaAhQU/oZLb0BFZWkYpPhqguwjxM2BfY
DHJgdhrnDUUL+xs1nEE392CfyL6zlGxvNduRF/bqM/XpXKCmn+yQqYxBdvK5B/owSBBu9kfjbwNu
Cigjyo2VEB2iIKXnyTAg7TQMd5Z5YEx5YARTyIkp+bn65pm9gTPrlhSCy3P4jqN0+5ZrOjDm0SBu
psX++yhSdqPPrdcEksgCn10CukP99yEIQDSPQ1etLErdc8/1ezbuE1bZ3r1FmCm/8T/NlkjW56bu
Is5Ku8LpB78HzOYaYjEhbJZKdG/yx/cHR8GM+ikan3JdcbSTvWIVV7RnbuvkIjOGR8Bg5F8V2vCA
VO3pyU0Hii1jBUbvy5UJIzJ5ovX47cuVC1eR2Oft0+eYBKBu+zZjHYTw0aZuZdrkWJ1JCCOzd4JW
OpwhMa7KDHSdzCbXozU3Dr8L3gzFFipW1xYkXjUAN6SkuT3Y2ArWpzfxR4I3z/xLO3ZcyATC7F9Z
XnWVkLpZauZnsjPCmktf5qO64BvKGOLpe9OgDFKjbpgjVgP6pV1dx7c9WCjp4XRb2eYCjEKaqg74
dwSzKn1DPNXEBy/Oy7FCPtobOGJlckFGE6/B3rn3KQC/iH9jRhrGTTvSBU6CC7UihijgZL0Dg1i0
VT3btjA6wTcfbKxIUYcHUFgxNkOZILQHCh/A1997d6sAXmZhfZgCdgDuAHf1WsvznFKAp4Ly0lN/
+UM/CtT68Kx6bcYOSfmROhuWmeE7j7J+gwzQ0a/rWo69hGZQj/CwfzvFC21ZUGP8c6Pq7wtOfHlq
V6sUdqh8DX6hYwjGHmGc/cx/Sc/9eHcvv+f+EKfHyUYWsDnuQEH/2sxXtcQY83MFU83bF2YOxhsO
8unfW61m/FKC24jQMxxAS2cNp6zMeK4KYz6My4D5RaUBkZ0oIpQ6RGT31ns+YKDq4PHSKYX9jJwt
dEk0NhW6A+wBMlq3kdh4CsmBvdk7N42Rudks1cfwp0MigFHnM8CfI5h/6ch/XM/PnwrmSgzeqbT0
tIoU1EoZcH/aI4j5e4WI8gbM2pGxzsfR0Fr8nTQGxoAzNrGuR5OlnQF6+of2lfJ0Q9uRrFH5LWN1
50kWbLMZ6+05dfsglUIooyOiHbJyPXig/aZYC7mpvHywicwD91Ah4xkwrauGLfIr/rXCguTqOGrN
MQ+06CNPJGO7sDV75jgUudEb02KOk54tOpmkDIwG5mBOrHUsTp9/OF+fys1ANJEvfHwSmx4rtkoY
pAE6w8lYZn+DrN/lSiGJlbrlBturYqArFnGOuq96/XmhEbA2n47M5Fx3NvlNaj/mkP2oq2QLoi5F
B/LnnTbmxeBef7A9gDpJjCFPGUOlurNz6sVlCpy4ezbXWIb/LcdrGdUasG8USDAznqQupvES3Tqd
YhYzojG/auzcIMYppjFtUCZXzOmM6h7nLqyYeRNLuR+g2niTdrBduKXPY/FJW4xHZf/E0kqALanW
a658u2/w6ouSDP7XzpPbsvpAcvc5XCf9qzOBp1i32yLXeGVe1FmVjrNYHYkcRTNhF2kHktYZMMAf
So90Ziv88b1RXbXVRBwHub+FPNBYTgVshn2n4CJzz/u8n2a0TBRXybqGrYVvsmGcC3reVSVDOnXu
khP9SgvxS97WczazEeuPlGTNRL2RFhCzRBM+J4RgUgrTPMM5jugZKcpiTThW+Y3N0vYg6n3P93lg
38c+DZRlWTKg1G+W4K2AM8+mv+wjLIL8ODnOhiDLpTH+HxGe5BQgvGcBaRMC7uH0uhTRZFk8KmGg
cZmDlMzP8Me+z4yjPK7/6rX75VJW0AD0+W5ZAfykDgRkiWYopFcE//E0aCJIEnWcEg0vLr6s5WPt
2VhksL10x7lT8hCSjcobFgcyRxPJdZQjjrZBy7+9vulnnr8gEnlb8CTA8s1k9dvakg8zgZezxMl4
YGe+oIhTBZhz0CToDsg2Q7zpTgmf35sjyfv8iWdxPkEvxVe1Ed7dtT06NrBKAeyl/XPQju3Zs1I2
Z5Omp9/iq9gMSIeAB7DTJJ6qyX8oXL9fG7qIG+uaN6gtQn5fz6zQ18Sn6ZZERdsXipytgukzk9dZ
W8z+EOq+4T4h6+rg1XU0yXbygSW11XpRGPIvepGAaxDzq4aItSNEiDD5/N9fTA+7M8zsOYcCBBQG
0m53zuzsfoazwhcaslZdg6TVvj+/zUDuj9+cL/UWgUVRH8LG+vBI4eOkfOSwEI3Ik/lrO8v5LrOb
1282B0kPQEOrErKrDO/deBudL600sG8iuJfFCN9/UFtLOmr4amuAkF4JjKo0x9oDlFp7kz56wj/p
3NA6rD0bjPLrXiUaY5koqZA8wkuP43xF8RlTFiRK2ZAb+QK8F6qyJuYmUuSUpALg8fXOjq/m9KB2
rrZEMte3HyjtRAh4/eWHNn5oTg4oe5X9l1OzO5i6bM4YOn4PAYRyeZVjU/FSF4sNkMaXPhe7yJor
Mqdq0rFcZD2uZ4AKp1GoNu56bnCMhV1Agu59DPWExv5ctnIUaF8TMRqPc92PaZ1h0TbGoK2zT/cz
B4iW/zHMkJtRY2UeHhQpzqjqlqJcp4HZv8hRWtZYL6jI/TpoB3VwiSDKjyGl2iBoTlkFBfHf6ArP
+zz2Qza2DQui0Jouyk7GCBA5mm0vXDzE5+1nCcFBptcrBbf8NzytLEk0YQfyRBYZ00XIkOQHUtHh
2PG20RC/x87AyjULxaUv2ghLFofnZdnmNKskz8QLubHE0Mrb+gfPbknrCMy1IBVWdQcIMaTh9SfP
OLMzw1+HbNH2NCqjkQvtKBgtSHb/t1eMMQeRfy6zeTtj8HQU/nW5H0oKB/n3a6sffFecC+DqDpqD
9QKzG753BhxjP7jI+QHOYUVbThMAnDFRfB7Khcz+9w/O24EbdJtbwr2T3LbY0H5mc2rQifLbz8QG
9wbRe1P060fGYM3+E3lvz9I3OJalkJfMcqOGsE0O8Xf54V46Gr31XlZb2Jck1VG9soOJ3vSkn+1J
VqVvqmS+cOMcvfMlIsDSJl5G3w5743JsvTdENueFqrANoCf3KiRBnTTaxlTOgcd9w66PLeHyFeMG
IULFuCcN1w4oNSokAE96Vh5i8hz7fiwOgW8JSybqjGS8FTNW6EA5Zs9qBvZBiDum8tccFHnJKWvA
EG68yE2ljfk3bmG2r3mKTUfMkIXhpPvaPf3zymfSQ0XOmtb8g5qt3ba8Ucoes/0oM2WKkbTAASg4
y73Bprw0A9txHJmS5NpqjQgNDQIkWW3hbkV8888Y19c/agcAAlS5g+R2ExpROtYG+fQhRSj9+DN5
XtJZKbhS4C+AO2u0pnKunDmDh6xSKzPgGYb0zzGJCXBhHxeL3VUmeL4Lwb4VowTC2qfyY76lS+/E
25vTasZOntdRHcy7vmagsx9Na3XcUtgqwZvx7n//B+LaUBduvoY9Dqov/eAXvDWr87aLa5ODK6pd
6Oc1QxmmP91Xr2HzBhPcnMMg6U+EP0tsFR1oWYafv2y36aTgRlvLb0RHxGTY9a0V+fIorIoY6exs
jCvU+SqW9Y4xnd8zB9BNv/AxKTbbMiSYeQdXEGeUGdJTKa/O2alH90buisZhj/X0bKIYUt7xeHwy
Stoj1fQmiWkRlyVB3lib29bxcOLNokJyphTzFbJUPHgty4yux/wnbb5fZrxjyfZmW7IjR0UjHzFg
UtbuigyQeMcBQU8j1dGt12eWHsdssXuWGJfwBe3xoBdGNFWfjg0W00mLBYWNDOmRj4ca8LVqcMOe
pC0wi6/CBb8TJGSHLDKr3cu4z4rOBetDrQkTAk4IaLscIZAROqrNZmPH/rIgxelr6hZQsfhfnRTp
7Rg5Js+Txr41dQL5j3FIbG1grpMvN82JhvdykVvr/aNIUGqkNuqjxRC1AAH9q5yF+IqNacijsIoY
TQRyfv41+Wst3cM7HL+sKgg/1xXCmZEsP+6yweKJcTTF1Yo6scZ+ACxkJfQkOVvjC6HMb9oSgvjG
zK3efNkN4gmFIRyNRDaM/vw1KEKz2Zd2TLwvm3eale+38/0EQK3gVwfoeK2LmYl5WtpdNTuVdk25
IljgMiG6qAjmU29ItExtae2zEekayMRTz+D6Qddsqj3EN2PjfFmOvoTHNnT+LWHU49MdI6wEXfR4
mij0p2r75xsR8lLVUE4a10bYqj0s+8dsr1TuxiQj09TBrjl/iDtr5REHVQ+tXoAk/1C4OXjHshUr
WiwK91muUyCKg3ZQ9TrwqAeWGeVWFCbpdkr4dV194aU6yocZ6EChCHQvr83l3tnj5tt7Y0Z6mpkC
cOny562w7tWibSg3e4NVHIcG2Q6CA57Sd+NZjxFqCaFL1W9E1KjVidNLoiLAWYbkTACHWDCY/PpZ
yWx8aQuyRs4ngC7TMTyNSxImp5WvVpfAsttx8t6NpDBJbp9hL51UZ7/HTmSJhprNg/MftaA9GH4m
lWdiQUoFKdOntm5WLWO4rb3953LlbuvyLYQb5vRmE1yqTbOfVmy+leBD4MDf2TUeuJb9t88aj4KW
zv2tv/PiVQz8MbeZhkpqSI0Osx1AVD+XCqySA3oFwWQFlz96PjANMw/jHg2GuR0b71tTq7/Luvnw
GfIQRUNBwZG9AviuzEv7JdqVcC6Qs8kMpeEf6t8DleDtYXRniy7ZN8uEvfonGK1FuNnMtFmZZTtc
cEjfl6SBsohJQ4BvxvP6k0OJGJso34/MGXd8m0beV3+nG/wAXInvG0KaoioIc86F1hlmMpaAiFVW
lWSGjaoCo7eH4supOWWibYTrf7Esg6pNkPewW7rG9QCAJnCYcdukB0qPEEyXvgai+zBM3CWs3vNU
pyz9phr86VjL0vXpT8ctJ3W8YbbcErQ+CUxj2TqMNtuf+fwxz/eNpHoeNKm6JbmDAY7qUet9aYxO
f7n8M0A/yph6Sqqhgc05Mt+8vG4br0193jwxLLF6JNAc2xintRyeS+xv7MlmCOTYhXyBnoixRgz+
qpo1cri2ckQmOKo9sR6AGLwugvwc5MSYelLgkLsf5naGiN/3HZ1ncbZKK9JY9qYsnHo1UvA5D0fa
GfCdvtmJi4oUaoFD/cenIn9Yccf2/5d8E59IuE90nfQHeoRmbtJwCKRdwkLFOyjyUueMXUQlRggk
7nSEiE9Ddxh+tryk14FtNLJw2qRxrmdpKEiO8U8p3Z7D7MzAHlBVTJVdkTD9Ck3xYb8+lkW4zLcc
xqFqu2ERpS0K647aEtMsYDZ3E5XQPf5f6Y51H3mMUTnEk9CeWXu+7Yy7M6WDez87HMhwLJZqDWAi
N/bxohII8U3z31BLOaI4fHt/rQJ+eDg3RcQfOr0ilxOPR4bVNk7GDQNXoxbri06IZqmZ2Cai+YIY
xg6OrtfiJ2yUV297RMTfqjdr4oFW2vXn99cuX9KX0NVLvecAIfw0Vy2RVkT28IuGm/JWowwI4nP1
1eoNn/DMLwfFCAsEtZf7cZkQi2GE3MH0w8gBy0KfZcHFjFNNxFWiCxTdnKphrGJ7uuTut3MXVR2m
VYwPWjWnXZvb6MdUbWvskq5lzUEJ+RHLJCpmcDxMEXihMnsBK3P9RfOim5UHQI1zQZymncQ/wNLg
nrK7OaSpd7sfFXL94t602k7xLhWnHqItHaZkG4IpD52h6V0NOgtnqAaWmG0fqgZ7iC0PspYzXsIT
mEi2RqCiVW1p657WVyJkYxyrxfn/YWikFp3C4N4FuH6IhmiuTgIpWQ7lT/hxLpfGbABgyAy3WSGs
le75pmHjdms2CXFQzUzoa+AfR0vqBIp4KFBGMBM09FpOS5O3eISLz2aa2Njl5hrKYKGO+msERSIY
OSpB38ppIhNzKByntAtKvUNdl6IWFLtOFXQoD7VSGLBvl8Ez37ENhpxA6wTtO3W8Cjk46ZdYcbcW
zn9kpb3+9+4nYNwTUASkj4W/FKJUsNcY8smCO8Kj4FGp0rjckyq5BivdXjoFEttW6UE6tru5fOlt
z8t6FNEDRGXYmda10BFKjE4kUWe7Kpv8CM149g9NSQXA/7a1Hhrca1n6x94E89hXN2tQlH2nSibz
Ox/gXGHSsEFlHLuOU3GhNH05II85P/vL5hpD8P1mDgxlPtw1bkwSsWUJnDdMaq0PYp2YFVNofP/S
WXJRpyJtWmxf6d6wwJ9+50wl0QcqAIjWfQrfxDCnr7KHwp9FeyNKBzCyj/ZwGPhFeHOfu2Lg8bHA
MP7hMUmm9d6avPejNq5I2EZe3Y8ehFpRlwwo2UV2c4mZ3/nyEz73nafQ3Woi7PRU7E4FvRcBP4cZ
hUj7fDCrJ68QyXPNsjPpHPv3kOYAG30VeTmRrSI7HMCRpU7nTt9bkgoHBLpCqin4hFsdT3weVEue
lNp0tkOrQlCerdeQVRGo54QPIzklehf5kbZAqzAmngPkYVW26HkrwJ+D4Pjbfxs39ByCPZwAtXDP
M6/iLGU4FlZ5ulfI9dwdNsAw1y9l5/rEmsDMalXjtdRzCV7Ha7vqx22H6wJCDwaHI0gd0eE3pHwe
vHorCEXnkEjaRL8KsH2tJAQ8wGr0XluJdQZJmtcSj7I1jRXK7Z+sKNsLwrHfDEd/a8eSGOaRHxCz
0tnTTu4ACmswz6sSc9PqI22Tt5P6H6a6c1C4mITxEPJ6W+fVLBfURFM21jEX8Bsnauc6oLKrcPRd
uP0NrnHhsox1GPWs6ZcAcd3o9hIrKgODKmDjEgCLmlHp6CQT8WWsU8Ep/MZf6LsUexKijPeNvYtE
52nxwQjZB2V5ROiYBfUkedq4PiTiMHHG01mH9Hvjq2bfvau/C29k87tGBb8fetn/8+h/azpaTntL
8M/raiMN0mQRUO7DX7/3VxDV4/S0Eq5Z6VSFVnHVmUFP78iLETK3smXbXty3XPYzwOsyjQQiY41E
iLzPfw0RDdOltClcX6Gyx+k77XoMwrvZF6tkuscXZtLipQMkZSYcgt0HZvhxanVEJQnE8iy0wwfY
Tf1giqNy0lXzQQSzQtM3YVmdzkJyVNUUKup434QqrQAcIBJIPfEbGuVu+rdgivKEAANsjnaF43aG
7/09CQcp+5wFTh+6NlgXnHwTsKR7M/ylpix21p+xIjMIhtZG2Syu7zLD28TIilgIHeAC8h0Hsm7+
zZFP2Vf859p7mfuz+UYQTVe3JWcsf8CAsV885RnIhLf71iIpSvu1aE0O8JQet2KLXfiOnhPaVdkz
WB36IRS9ALhtmmQPO90AeKgNKw1RcFnOFlDZW8OgRXApgWuYDuHzg7vSDtPLNGy3pAK00YHj6kdp
bcn2LZ0XQqooWSJ7aJteNxU8Xf8mXuFwklC8qI1zeoIzPFEWbuxhUR+/Wp2SsjmYE6AIc8ZoM0eD
jl92SJhINFYPme0JYsYb+BMDASKdQGSErHvtj2EnPxQMomV0vbAEXwxsMEWyOEq3gAfiXCaep7F1
Wdc/2yt444TF5lnZtpRrBDyO7K776CZWuG2SU3+93QBdYDJTGLQhWkp4LMrKqFxlIypdBbARDe1f
Xee/qkIxHmL7aNrlufzdFygv8NYnt+LzcebCBfwSQr1Z+rh6MBPATmIH5Ye64+9KQDAqNkty1ocC
9Dm64DiHBRBmk4DRbRCw9WzslIIPu4DjXtiMVNWf51uxQpcE7Sd5NLvIM/QFM5CKq+PkoIVcDdnh
az1VNIeu8gU5CmqUoiv+pOXVb8pUpGAxvVr/SLb+a0uj8A9RQIkk9YpIeZPfaQVdfMKKXvXAikg6
AZL1UNPZ8LwKCYU41D63BiCs+XW8bT0Xib4PYcJPdCAt5gVcYAV196Tv9OzghZNqIDqd8Gpa/t91
etbkGayUV7ORXDWABvQpnkJZAAy7OmSbbyyM40Mle2Y+Pooz/vbaxudhLdlXYNugZkCnE7quo9uB
X2QwmdI6f5ZQvogFfhLUQnIJ3KUGLS69ATGMf1/aJKNKJexGs+xenHOQUQ/pG0nJiZTpFggEawag
u6av405TnH8IxVIlzqbpFqgOzYqHVSn1dgwh7ENwUhPzykZ1c77vGvBy4yFcGnIl9+9267wZqzai
6ROWvTlulWt10yq/VbrYFWaWEfinOOskVUWFXbCeHmQJ1coZ1xVsfm4rvFCD3NDTeUEllQFtRRof
KzratXN/E81rP9dJp0/h0HJxVY1oGN/4aZMxrflehA2fStzdqruhTwzv5F1RITxpcDNEW7TFqcJr
P/shm2cfVkPitaFPke1yP2fTFy5KgXfjsVmAdHHVgNKULLjQB4GXDw1dVo/EgzBcy+iaIMgiXS0P
XS+RB7BH5csqfB2yW38XiJF2UqVurAkBnZaHLE4Y8AbP5+40vuGpnck5+csNY17hxEv9WYBh1lVi
OMiHlzIxPFS3xZO8XiYhdcNTKfdx0g4UK4UTcUPQ/G+1Xk4tdSvDG/9qToTSx2EgdfjjiYj9vhEC
NxLt4lkRSfX8vGS8TpsyjOZEhjJI+O1x+AvCANEfxPVotoXrSEIowT4QHCLYNwb3dBI+wVQ94/1j
qyF8VFQp/aKYzUav38fwMRX2lXqKtooJqg0kAEx+0Gc9WW1expiaCUx/LFtHU6YUun7qDTVTQ/4j
w3g/UjPnxa7w4RLgzQ7fTIw8HxzFoF5FcCU3hqfbeg7NkE54hdR16s1uGjw9/kGUpWJYTVtnGDuf
e3yKzwDn9FRyyrHuUiOGgUapMQK+bviQNApWp0roF25aRwb7yWr+K/Cj9vyqrpzigT6tjdL++MuF
SdMjrnPTuoE0x7iH5EhP9d2m56EFbrmCZV1i77SWA8jJLwE6Mo1XvwSmUuE6JUieBIyRhh4ci0BL
3BSLvZrP2aX1w2AveaZV2oUQlLUxauZrL+o7TSgD+OhYvYtTUUs5g97C/2A3oNnCA+xLamPzGAij
vsi2CUgCuRuQy43ik9BHEopRZMNjKfuT0LEdzgwSAxJLCqQ3Zdi4p9PRtxTmCkpqxs5O3H8fYKN3
G3rRU7K/1wibZEYuQJ7YIX+qU8yefBUNpRGcj0K57Iv9sjiuVqv9nPQX8/A7DgJ7GhOe+eTHlEF5
CwZ6t4JUuZrr+/mz3h0rnfLbENsBY04JcOVGpI/40vdw7+RNGrTSml0XUWlmkox2ZcuH3iUFq+Hh
P53fTaWgZX4pWWU1Ip2wXWFMOMtozq0+5HOTXVgsP2h2SnJIVYJnK1ne45o2M9H5PbAf6alcuBld
LuAei7qAYT+6Oe0l8JrR5caxeRf2psNYTpt7ycXJ4Bua9J1d6JdS9cg9aucuvsiakp0bi2xii7jN
l0hpIKADuL3azRYmSiV+ZxuoceYcrLKYI+PhhHgadqc3HVaUgwvvU8zUnhNCIuA7Jus6CcbCYwP1
Zylk5ybS1AnSuldGfMU2hKFV5c1FoTMAeZUTZUrJVXXtPb05y+pjTbIRHEmrPFOOrF+/K0u51lka
wqGcZ6L/W18hSQ6BO6FAL4OrszVcvuidpo3gHJtnePI3MTGpy4GvoAdbKDdZjNMsJbO1Zb0hy5Yk
xIBikAbkq/JA5HIr/zxFrKwiU7/FT1wo0656vO99Pg2Lfrzkc9DXiCXIWTVOznUVFfWj8fFcUIjC
UsMQQwAD+gBKx65Le1diPAua8inYBpiZEDI0Pji/h/+weKay3S+8rVk82V2XU06yhB1ErGKNPmM0
NIok7DKfNcRIit6D+dta3Jwde450KywY65qfKsvby5Sdv1C57Ma/P8V48zIt/MvzqtrhrLoqWTtf
KbKfMQDUlkrFSAmAIAwWlzkUJB3ryNOwznL8W+61/MA6tfOCkyS4ziCGZYs4b5/mzu9fIpQCVVy9
ClVD8P7z9GkgTTd5nRC4L3+f3co2ug09jzV4rp4HyJgKK/UcpLvGqK490KyOJLOzDya588h+EE1D
Ortg2jRU8qbViLFT00x+RBdQVuzEPJ27SMsWqRwJscj2pxNzi0UR0aPpczeYxKcGmVkT6FosyN5/
uISF0sMesSUu9b0RUyibZaPjEL/kBljslcrOSHXzXm3muvgg44DNEmI2bEt87PzwE8N9plYz9Chp
tT859pvp0AgAHS6J4Q9OxgDSYcrTKNnzKMEizq0+OoPQ7u/TtW74s+D7jonYu02bctx9RlO5woVa
r1YU5UFGANyIdtZqa1Tu31lEZ+qLkhMYhRvXdLgEl6RaQgTBJa+DKzWSXoQ4nwWItZwfVuuRfLVG
83VxeUn/TMG6JNN887/Qw+qnV0o5D6neK5ofzpVgxNKaMcXkf5OcZsLeotmJOwB4PaGqWVip8ifB
CQcFgmAO2QBmdXtIdCJUtYm03TSzShAovfGmnl7mQQJJbYUVrC5tODnjTYTjjoRVf8bRCyPiY9Gg
7K0WIGa0IHvnYje/qNMQa/KWhVduHHyccfeqDhx1huWvTWj/7T8Yaatua/aMR9nsS7WCRinVUPCT
1bNtIpxOPX9VgcNY1wWWn27yd1arOJAq32RJWtGpAneHeJJoyQqG6e5AYJeiAKdWuU0SObYAFWG4
oTd5ir8Lpdwlk/OmE//1BCbUhlgUrwJ4kcDGNqmt9iF70IFLJSuss43+0VsML0W8cDTpa6Xm7k+T
KVrjcfnhkQh3B4FN7mFsQjwZFpo8bJ3Bs8qe705jGlTLLaLgvSB1W4Y/s8EHfS4a4FBFKtEjKDjC
a5Kj7cd38Dd3QpjUJLRuEi8BnOhQX7fkPqGgWG+R4RSh5Aar19ZHB2GH5ewQFN4XDbBruvVhvb95
qx9se6ZhmYRQp6i3EUmmXtDfX1E3vezhsCykOkzZlrFw4cYi4dq5B9fHnUebwahVgy6tzewbP6WG
6+/kQOk8UqQQmq6SVV9UJCMf3RF6jZIwvEcyhjkpT69FK1QrGdsMLbxLQ/nqAi2OLSza40l/yF5o
WnnuhrmQVIBCHcGDY3DWMNwclkfr+TXAn7A2UE9uANO6aXisniOMu6gc7bcQQ/o3XX0OdoSWGuxR
YWxpFllDls83m7Tkp76sz7BAUpYzcfewi6forFCyxYV/lMihoMToW+Qq2yg8tcBU2E/zQQXX8QnG
tEVeogXyXjNLfAWY2Jx+JcVF6r+qWi0Rf+sP3EfSp84bqxJ5tOfYIoQCk2rc5M9eAmraE8KqwP16
ebymjtL3Z/odYlYmvSJRvcR/FI9ZqyfkLAfApoBUE50o0iboGy+I3fRUeLWXFEs5KHmsOdSfjvYA
1o9MEfwt2CCxTfPXTnJ7o4R04qITjWE/YNYy3/NwmrhMgGqW/WRlbmtu240xSopMWdH33ZjPvZyi
6RvLsJ0ULLqpKiC6tHQ1imwEL+lWQpOVEvMxw1kmJZWu1EL6pZCq17ylFQoE9f6TAbV8vwTSo0Nv
EG7KvXD186PQ4Mmgh0cgQio5w+eCo2paIhuoYuiuP+CoZpEigqDJ6iwYNuYdP9kTIzwtlZgPXzVl
VNzgL8FvRTXwUnm8BWXtVmrRXfZZc0BDjyreE7oAv4bEjCHPMs1gvZGC2sCniQmYQcA1kmVzffAF
M/QC4ErOC302/Ed1SpEIjJ9RCP8mamQRlEDAO3wSnJbOgZWEAk1y1Ur6BNL8ZuvEFVrcA9ooQP0e
jzxDHeDVopIZcyIT2Tp61/3HsDgFkkfc3rk0fTncs26DjQcACN+ZAsJoIXwVXtTFPFfZuWxtpkHz
ZcETkq7HkoxwUEuz8Ai6rce3WKndPW/nZ80xihVu/o27kig/qUh95mcSBAXpEDvCIL0bm4MwAjDH
2aYMBCMVfweIhmPKGsK7iAjH6PhLhSgdJs8LRSk8ZwphZm352PgVB/jMoJu0NOEBWOoyCQr+0SF6
gQnj2Rw7NwLkMi3ssQ3bFiUCTChjSdOoSpVkZvZEMZVNS1a3TMXv2xtiefsTZ/Upp1Zb8evzgdMC
VR+NIR5r69bLGvfDC1qRoKdAdFqTc2FAnNjdgDC55uS9ulI7BfLLC7sPsViZPwk1nilNPqolODkR
lCYBT8Kb3y7o2wUIq2NWEL859st/DlpnC6t4hvVaolJ0W8KUG9elES5EnUfmyCzKO2xexS5W13PV
BmfSB2GT+vvNE4DQDMIyrx01lFCMTo2GZBw44kARYpZJeYoxhS2nQf34Ggia4n+QdK8VQmoV64Hq
ubt5qc84MEZK9yBnKOsd2QVLM5jIXkPSidZPMg/E7LzIRuP4i/iamF4DeEz1OGhWYRpbVSE+VHaB
7AIckZQDeB1yoJHZsIm0UygBWueX3hxmgNqPt8oJwMJZrQswZUuauwUywNwGK7kruNsG/aGDkz1p
MYbRayNPkScNPmsC2k2jD1zdepyLHW4f//OeyMvhcxpcYu9qeCuCsLnHqVsocn9gvr/WypA7xOrl
IWlCDsE/2OU7Yq500Yp9FDsXZVZwrOXjZhm0oOgu8QZ4StMrE8x4qhUdhoUlEyL973/hY0rNTaok
SDOtDFrLP48kARk+xuMohb0Jzt/9Gniohu0WUg5V3dH3aE6jY+x1wQO3dvCtGSHzg2sFQm4goVD9
ounBLvauPLs51mXbsIZUfxmEPcX3tbVgpvmq88fak0IFCrtsCYZ2Bc+jz0sgxD2izbEM1aUgCRag
YODC0vyOyzw6xk4VClfqGEBvZRbffx4Z33KuY7Yrv01vVVcrVA0101t4IbHBlGGV1SFUxttl/YvC
7GLcF2jsaatzpOX4MXZtHTjsTFH0WpnknSaYaBaK/Chq5sx76RBr0dt0uyYuMlEtd41bt0upXWpn
fk5mPR2MssxnxdLyBCLca2I3xY64bwW1j++zKdkahDY1FKHRmCq8Jng/FTKJ1kO2NQ+HMIeOx2SY
cUK6Hn/GxSpmwFekzZpNPydIl8dSEDss68UJGWF289J0tZe1w+K7P7Yp//RKQJ+19s6e+D3cfmT9
YEWqnhknuyDj5ECFiI50JEe4RjknBierEnBAGvYSiEKskwAn5cImDgILKhQlOzmqMg7c2/4KAe7+
noDVdIaskMP9UzsComExVufgu5+9azmcYiRDtFoVTzl3ULKV2TbakXrv75Ol2mFPmw2I6TC/JTU5
odHPWQEr5nSJiQvkHo7x0w355jL4ZIBeX8hnXrXwVcWHiGou2mqphFUPHUtw/WSzBGwbDral2C6p
fLw/+Ago29ytNDDttZ52Mfu72WBbPkQjIc6L4E8HOYDkKDfFn4WxC9K6s+KGs2VlqeP7yB36CG99
pxADgqAfjuh3KlOlAmbZn/nty8amJIXkRVVwkL2WbThfZRIVdzze2tikbo5rQWMEPcBQ+zJv5+3Q
r8CtdhJoJ25C+JO6yQIvIazDbVzzYIVCmx/8nA/wYiFsFkT7RK98EbEYw8gsA7YqpY5Bt1DTwlrq
i2kodsTcYp5zY945ZHnNx4BZdUUgF85mcE71pGlrWQI8qCBx1MZMl2yNWzqNsP/jS2qRIOQj6xGX
Hf8Zf00Lb0qzp4TkecWbZEkDPjl/ldzylFwEKxaefX1Xv1RyOl44APx3fYthE3YCznLxFXQ2srzu
kX6xJiAnG6TTD9m/LHL6puJwq8SISkvoJoBQlwQzrlHAXi5NM8UmaXKrhTa4C6K9XWJayB7or+OR
xzhLPaJq3LjCLFmM87uJVI2FZ5lCsCR4lblBHqZfyRKjEFfaTrs56tWV083pfiDls6QjmOXzXdCf
DBpaRPBZ8Bb1/gKOM07cpxi7Gvzacxk8MY+0eTRnUTTptM7Ix+RRgKKH6pt67bFXYfaXNPiaE2uz
0pOo+z4zAL00mYK0IY2ez90+b7IMtm+cIYrcumeAqXzOI5n1dHfWML0o+dbAgyczp0G6B61tNGdm
+mfey/qBRcpaunaRhk8J24ZOh25QvkKJKbBZR2MPMAHvJprhUl6f0w4H26VhdrOb2KRwsjykFuUE
u2muG6f1ziNB54YjoJth6Bck+jHS0aRwcebTYlESSuFmB7UoROFIQOqVeGKOloKArQrZxjGl8rrN
+t3dK308yk92E2MGj2YfEvaFkBKNWxsQOm9TwONFxfxbQByCsvKcC8dVENoY4sUHjfTPQcgSA15d
vaeK25nXKlgaqxQfsf+LceB7MB9ZPYJ+fxiWYZR3pydgNK2oAjwrUx64BghKWJ9U12S8lr3Tx4sY
kzfweDcqOlguX2TR6PZklWJmEBDoTKlj95nIawDimMWJpuHHrc713RJ5ZNumC4ddaZXVenM/z1iv
RzbQ2oWruSoGhqfjkXJP8AMQTY/xVU09QHgKeaWI+BpHShO249ZdCfK6Ofc5ipElJY0ywkIxiaol
6T6kATmLkn4xDMBCObIeEbxbzHyegFM+tHg/dRdY+1fg7c/Z5b2JIWYle4bH3yI6wAaUrItdEij6
gVs9IrlW3D29db9tOhXkteYi1rOTwfB1suJ3oLvvY+l4ovQAWNRXEg7+CHmnO5m0Cso/+GKyh6eI
Ho5aR0wfHPT5OKjuyBVQwrLbTSD6Hdh9gJdW2H4VPdDy49NjApxH0nCMKT6JImwMHEyhIBqHeKEf
bplbFFtCzEzWzgktlSuYdIW661idFAAu3XL7VhmLHVh8ggDT6gt+bmx8gIi/XANTHl+EuFU+cXn+
vxEGfJFLBVgVlgbJ/pWt3HlRL3+QMYokonLegHJ9iRwk4NOoWQ2mFBMeOdp/B+JvyEA0siypa514
hnG8c9YWWfcokFS68/hlosOEJnXPq5+ic2pdPuMSv8SSGvNvpiWt7hSFJSW/nbulqoKoDYbA+RE4
u6Qypy9dg0hHp77T9Tp0QhK3TNzWkaJqhtVd5iC6J8Y7EDeyRiU7NdTtLrDPbCPubNqgPZzV/Fsf
WNqg+FSok1C3EsOHnBzaf5OZm+UjcFdGXxR0gv7oBk6xxfVNf+Pards33ARfQCZYtrOh4KF7OKNR
IfNHQV3mwrhWwkypGMpS4VyH3y7jtAXx4g9LzziD47PBkcTwHJHU/YIKel9EKIWId/TUe68+PR9C
Yp9OGnVZI52/M2OBes5SoGb7iN62AFmW3Gv0QYEWOtdMPw9Pd4k9YuluiUj9NeEwUTpMui/BBwOh
DuNT4KYZZ9xdPrBd81WU+/fC3d7V8pS+4T9IUNJMRHKKy8Fu2UvO1hM2hNKeJSVkb+Ww+xc2Cjha
3PUtzYfdD16MoLnn1SrGNVz9PNXaid1yg/93jPPk8aP+lpMQedKr8z0/gpZeEXIikXB4PuuV39S1
JP7KNLYpyg5iZIVYhCNDt5fgmE5GD8tm6XZqOpSvam1vbDRMJO6h0uNl5piYslKoq1efd8aGeRRU
/c0VmGRKBsHuDmIsjA+c9as99uUP5d1AZNwUsZmp7NgGpCPTbL05l0tB1wRI+G71gQlXpKm6nFZp
ki8XawQy3Dmqf4C8nJJZDAD8ZTw1HqXlSHmuwRhbdMSudB2C9FTV+hd+OiE3qGra/ToBM11iAtFC
WRcZQf2cgahNVW13pvkmcIvlF20vi33dNoUN/uBWick+xT3nj0KauIiPL9MnMVB/0adrJf7BRMf+
jqL2u1R7h0bP15UokXE7gj6YlzSIXPUFEy+tFwYAOKaaGKwdmF6hTHUureBo0OHlLxOwW+qmfL4q
L/8bMqI7y6KGKpqUWa15/LoMy0FHI7inqCOCLg1FSnACeyDqbhwRuaRBMlUMUAjPfNiWWfioPpEb
NfLknj/nwCxJypHRENIBzZOo49hZcHh17Jb/sIxLSyS7Qevb1S/wPe6h6vl2DRRdLDtM2scEqxtY
ybpbCkJ1+8iLe9DiRaYGv4A/4mDCRKI3s3oM5g9rWgba6io8zzdNfYZMffgHAmB2awAuybQkmOIU
l2BDmlYorfhW5yDpQYO8B/45Ts0EWhAjJ7Eq4ToHIh2OoIBg5o2Ci8XOD2oOWYUSn7WA2mPW4Kj8
bjDzFZOk4D4l13vUPOKV71ZsYUUS/rIYrUXUkxkAyRSm8p953YD/JHvyvoMPjwzG9BSoYp5L9Fqm
34V4k0iLFKEUR6uCvLXvW12Ss/evHMS85xH4kIkWBdnc7+3hfds/FRDdmXyr0+z6B+U4p3oFaKoD
vTrapompu+dX4jgWfAVxUg53mCZcovl0Oeo7lyLEiYKEW5VHaMmGXFOBu8GaNbPIlf9lAqAclDVS
wUnCtS+9mL3Jn4S0fwNbcRvxm3Eo059mXH2As1PNLHtrAlXv5pDT/e4FK9CHaXAe94Uvmsg104XI
UqLtnPPqbmqzUY3E/7iOxZlCNaLn9tCP1QwoS0YAcUOFYuLatYCuqS8XDby7HZZ2ptlWLA6tQlmW
ApDsayyG/Rh6CbrKwyJVcloeQPXlgudn8VFVo6JWSRd3kS2XPExmMJAK/vPoscEBoOHwzxLth+QF
OgUu1BSLtknCLvGBHja9NhqrP7Gzy24VyfqUHNsSMWz4LFQIcIHr7rEuozzJ+WiUt6XjWXVEt2mH
JjyjRorLuPvvnC0GBH+dPtBZz4nHAkitXa10iu699OjW/66SMqO0XyJCgW1sQtx/BeTcCq4pUSXp
xvxWpUD9S88/Pc7i3hAid/vXXKfw5bnbw2vFwJTBP9vyYCps5RhoWRp/fwrBWgmXsnbods2ftn08
JAsMhA/XulaDYfZNPv00B8Ut3Pb3t7QfQZCeSj/RSwh1Uf7TDfCi5GVF28wa4nyfanoK8khfcnBS
k8AW9mThq/FSUGv/jhpg+FExs7qn1u7Hf5U/7M9z4fA9b9qZ/O0vgm2IcQ7MLP86Jhb087o+OUvH
9l/LfGa1d1NexPT8SrAyB8kXKPXF4D2QHsOeWFwZirMNHAhT0C8FKUe5MqxZT4KFkEMG/H9Yeclq
4BDrgwRMI9GOuOSqXM2whXewsTE3oBVuusdW9mwMbvkFgORUQ/CswAXPuCFKPZQOikE0q+IGg2bL
/QZY6gJWy02BwFueM5oGaFBK+cpQKqg/mW1+RfcPs9yJbVT8KROR3CjD29zhvX8+QK2cSX69zeIt
rK++jnVnwlm3w40zBrq0vI3q/8OBQvFjwKI2klVU/44zep9QFL38nhvtEOgYZMJTMEIeu/tas9lp
itrzLnoii5jaei+cL3RK7CYYb3ro4gumgyESJoVQSvmZVYwhBMWDCnzdOLq9rCjYQy7PM2JiHCyZ
WILcrOBPRgpwySr3Kd0Cqe/k8IBbLeEy1vDtvn/ZTk2u7w7dMTS75SWl9q3O09BR4ieBOC7pDACd
51g3lb28x/QVSOULe/ExBNrkXFPO2O1P2Si73ld2Sf6ZfkOaECpGhF08RhPDhnSuepGDZAyZJWaT
fplbAFxEr/7vx009eF7iL56Mt80SFw8Ih8FquweguVcKe/avd1fC05CXmyc57C3R3JMa5q2Yg5aG
O5M5XyfIfiL9q3dE8I/Q6CZKwsH9A9tjkX3J9Tl3y0RhmxOlYEeWBesSl5e7zudRz0sXNxn0XEza
k5+L8zZnWGwlEIZ+alnWesz5+OUQiUVkK0cooC9xn77/qw10mnaoCZVcQZW63p8IXVhLLTlZ8A3b
QeTJA9azpf+RMZg4VVrHUY8mM2U7BN1gQJo6hoUEN1XpMLam/ZHJHWyNEufmyqsIy2i6jQvvpPu0
EYyTxwUCCaCcC26g1n4CKR00hKWYwPoRFICHf6kH5VY5XUNYRQTmMEz284pYRYmLSQdWBeigB6fD
Yqcr64Det1kFzGzw8snuxRQP/E6GK4xFt2gihclnnmBkikZkaD1fvT6mVTm/VM3vzcRyx0xZ4GBn
1HvJqo7aP5/jls0ziUlBMwuix6nxIIlNhnd1vC6t9URk7SG6nd5gr0CJUfmE47OQXcB2w73q2ZL4
PkxtSEKBhQrGyh0aNkVLtjBHrnTifE5IXFTRVzqkFWNkJf5gnH5cpPFOUb48M7/mi0MuaDy+El3y
2STR5z3NNgG7O5d+BlOrcSxCVqv01NXIf4OV8XE3QLfNuul6Ce4R/VFmqB702NfaJZKFQqc2sz2+
qkcu3BOYb0YJIwQtOTjh9fk+Nu03+n7eF71UZL9s6fk1yniCpyW00yMOfv+Qv8Q2uB15c8lkR1uE
frJsC0/c5tJCKTOwO3XiHjJnbMoS1+2QWH6wceZB/RYPUWQbKubQBg04RE1LnEVrpSOfpNeKUsdQ
FnZIlKmvaGbJ4gviw9udC33AyqbCGKU77ghzsQOzazqryFy9BjsFq3H9oZesFA8D2gQCCXb1pv/j
TNR6/n6ROrc/cqd9XBtucoRl6O8DHpev16qSmCrQhCP+F8i0isB0tWQl35qg3Z9zcMZY+zTS2SJU
4Grb+q7Y/Sc390LZaPDIt7xFzaEjg3s5a5JcIdfthT7EBJjGG9v8ZmwBklil4dyiy9rtV0+6GPVV
9uiCIa8x+8VzHxgSRnJes37dg2ROe+RPZK85IzC/S77actBngFinc4rIbz3sQzwKBlIj7kfrSC7J
w+25m5elHDQ/jk30DCj/FcBxzpIxH4vNTrsJACWZB8WYcQFASskh3sZZCoQ8WhAQSFFktBE1QGOg
8L5rk/diXQxdU2b6g4ggFQOxUd6QDYPS5kdvsWqyRPJ5m8Zd5q50UlSR6EU37qmB1fLTieQ1w9er
QXaSWXBkH2cor8iHxYrqdZP9Qc5wRv4Jf1cl/+LMFz6y4q6SYCwbj5MZUWHgqSAykHYHfey3rX53
W0h5Pv95/Dx2x/fyXl1gAfpL/g1kpPg2G3EyVlRF/x+hqLxSpGu1R6D6U2P7v0MNtrmlfOwSJIX9
ZkLoZYvSUGjH5TlEdMDdbUGM7qyX6LjkVXmC+sZFWux0uyfnWysjyZjViFGaUteOeByd17YdQ5hl
zFmES+x+lgOamTuCGycaW2yGqaqAVluH3EJ7c9dsDpl3Kbsx+THqdvMdmHil9iQ9QhyMRWsebovV
8eTmomQc2mhkJ4EDCW/jn+i053Ty84O+pWzvM1WJ9DMYkdC5GSMTUx1hdVkOEHb1vsT4/lMuP86h
ZOhGkkX7lVs5LLF4P+HsgTlUAHzLoMV1WRds6ypUBvL3Lr9YaQE/I7N99qXO8FmEp5WVbeQItJQv
ayNm/VwmzHUX/1+vV44AO/rriDcWg4DwiysDnwphm9vBNkyGFBeB1QLYuEcExDE5C9YUJTydnHH8
YotlNMAW4bTo7Lr9+8TgNWFcfz5vr8gQhU1v6aepEt3JQP2NlqdvDdstEe+18yoiALOvFVB1wHVG
wzj/1uH6uElaF2Oa+cGPyED7CwIHzhkiDnl/xzm4DtvxUCEyL224/BixOqllCyKq+EiUhTTAS3HQ
y+ei/czrIXeuQ09S+xyf4vpY4mUFRlb86tFq88qqBPubnuuzdi12e66AS9JQk92Z+/JTWFNAGI9Q
WTi6cOCvW9y0WcURMNoPRYJIjLzlA5m3JmGwVl77kBHClkdH9aW9GOPsUCzx6lsruXZr6V6WEgm5
ZbTnJTxDje+i7tu7KRoWD3+5shkmh6cEtuFooz3c0rXy3iiAuk2Uf5f0QStUDMhEnzgFeBUqrUhM
UvsxNOgekjNWDzUzu3wH8z+eZ9ZbclNKNiTGPWBnahudotoZvSIMCTLf72RVJZpjjIBmXbijQT80
Gzsd/touvUmr47hpo8RcnJ9meQrYCpgWlFz4M1jTvDZbnXax5iRsVza/gvvE7zS/LiQGjKqbyyDw
aRSN5XtsXlNzO5VVgtFuqeFyzykSJu0clBSChlH8mR1CvLRK+jNM0q3AXwf2a+jLTsFY9sKg1DPW
otyTzKlq55brYm/tCr6G/4n3w+Lj9wfqrBv+CNcUXBCgn5dFD/mF1H0gNBzYs0CzD0nA1H1h4wRk
0MUho73kMA4sIxKmk5WdlegD9zStXk+ciXm+wcbgJG792jsWZaTuPdfD4gsFidpxqpdcktCfvmry
2j4yqi40/D3hQVrNxxxofOhAYl6sNsevojYK+m3WwuWIv9Un0z8wY/kPtIFqo6BkQ7Zk+rS7xzy5
Y20LOW30WsPtHfzPRubDXj9wsAlQ/vwPuHptB/N7up5n4sCsgupziZ5L4UeM8N5Bq41VLDiaeDVS
gmvOX3uEbGfKxog9JMb1q5YPSqjEciGfdEw7ChwSkbdNvDFPctWRmdxEFOC3kmkN5Qha5cOD1KYz
ZUg9aj0YtaL7HOzjcIcoVHk9QKySJJIHjkrsQz5X3seeF7GuzFWVdFtsTO9gLICDAHJINJ9X1MhW
B+QrejR7A3TM6AuvsitBMSIahuMe9NpCpCiLow84fU+FYF7NooriZLBx6A0N/Y8p6CjVkrBhbUHx
/AvYuujIHXbrH/o1tFL4t+fDxMqXQKmV7MGl++yPB9damkCwL94bPGgeISIT2q+JmMJk2u5wrLsb
FBeQAaGhd06nCGUNc67taLhOyurQ2sf16MJpv3ZaQmfR6fKraLlCIKL64JY8RvUKApFArkJ+toTZ
XBQM80a1UihLoH+K7WArEP6Xa02mD5Zi3F1mKDr9vXOmLJjo6xvhsS/K2nGS7CgYsh682rX2pjNd
msmB8mEYaFGJmRfbYBJWKJwHBRyHNHPohbzEl5L7K9CkSG6v1HQOsFYiC/ykVllqAHWzuWzhF26d
kxk6YMQENP7a5L1kRfwaSp4JkJcZRvPbD4s3QR/Qd41MiexoJhFP6/lR3Q42tQ8838Vb1axk1FKX
c7avBfciSqsSX405JtPiWZrPPXBK2GsBMjgw20lpXl8CH+Efr2gzeOjUUCVaWSEtHn80ORJqkNNC
VoH9X03T/UsEsDhZlQryjYUpu3AWHiGN0WWEY25M1QF4+JvwThTujbgLXG2DZlrUqk+H3XMhRVdl
whSO0YKxeCY10786dp/6WK1VXKnx4NtbQinRscXH3sFuZwFFS9KbFAorTt48f+cVcAa6deBNEG8A
PPiWu0t6XGdNmG0dCa/17CR6nZPo0RWIVY7KjddhiLeDOqXcuK9+/+AZbQIymCMjhrHPfp1Sagkh
mYF1GG4nhSorxICZKazE+RfRarzLBul54D+9tHpg7kZLnbUWFzYxYrXcv3HfBCE8vCJ+tWmL0sGt
YE3Vgq72iTztAQUAMl0wKbSrxTDGZ6NHS/M1+PGe0usxrnodLSSD1nVWcI7xLTTdCBHTyVGbd7Cm
NYBEMpuaBtFOn9oq8Hc/sF8j3tSr5ZcLn7X5+qZfUP9zGdr+sF89fxjV+h8AKWgLYeC2zflQAQ0I
klWxeuic1oec6kd+VNOsvWgNNh46l8Y6c/tgtaVfrX5yoozxCotEJFS5vlEy+ZkmLVXy6CQgP9Ei
a0DunLbsJ2AmHNzft0HYzh72Fu+hKcqPTe5E1foSPzmZgtj5aCxpus59knAJjDwy5oSbJqN/ai3R
OurY3H+nkkOozcESnHggTZUL2BPSBeWh6Uw/8ZOSLvapI07kh+ibEUJnG3X9eTM+u8tun+qqmXx1
GGF+PoZU8q6RklVcnEsN//9jGGZ5nt9SXCQANGfSXT4M2JYHduruoV2/ERMH9owf1B7NrRt4UOOB
TgfgTMXi3IKLZ2vxkBq7mf2Ywo4AgI3KIXNADmh0KQESfOmE2NyapBJksfQk7ZiQhDG6+jze2IFO
aE0ELD1JdA+nRcBH7Zstl2I1xBDhKB/KrbuhH5EIdQOmNaNQuxd1O4/07RNVV7l+r4ZSb9u/J5EM
UGfAQAQLG/UfjrLyzN0gVccId+dCMWxyipI5q20y6G9AZ6Sbo4FKa54oKfQuqrtRdAat/TGkPmul
B3PMOWsnwAjGsYHKmZx2KU1iyHwdF2wKrPndTI0iVPM2YNaKzddLV7FFAaxB8cjyNk9I6gAREyQm
Tc2BCG8KJn+XVRfKZ7NJc76KFETogol2rU05ZaaJlBe1+Si965r10iIZCGXOcGnMgvwVZQ7CCiT0
zt4JGy5hq8YciKFKDvwXWJ8W70Gw+QrA0nhBpnN5UEsm6dgLjkeD9z//9K3vbojajAK6uu5G3idf
fOIUKgmK6Y8R2/uoR+U+VdUShZ01olY7oCXKNJWF2ebrIpD3y7DVtJG2Ro7xAev6QGGxwFu2yoHp
PhRQeQMzl3rHPeanvMpchrc3m54kdxi5eb4lW2vrwpqD8ezsK11H398nSFhG18voE44yEz3YNN1d
XiTdxu2tgaWc6gJ0kVS48Sqee7QIeYJAk6Hr7nntRmUephIZTadEXf26tXijDckLu4EoZt0ap0ee
rM+JcuqGh95/v39IQlOcsk/p3gk7aKfA5NxwemvsyZtGPTmLvlV+AlAWtx7Sb6QAK3nmW2bK2JBz
Eod1CpLiK3ohWE9E1yxL3gq59CO+OspLgmn2eH2OzV5sVAWVsMbJ+uljZexZspP8zxy0O+X9QH2Q
NcMhWUqsIoinR1g1HxVB/JUcY4RdwXmmDHt0IZ3PH2LkPV/KZzQMxMZpzunjoP5kIvG00z4QOn7U
5m2TCvd/cDFVIagaqAny9dcbZ4cFGyAW3w3lQ4ZEMjjBAp0u1d/K5ZaguvtDU5qq6r9OCdNTxhXf
7rDxa09SnDrOFme1u/dDF1WTxGu1jR56P9eT4jnlKwbn7blPgQnGdj+Nq0uvPXvIJ95FiIukmugT
rS9FDqIPEz2IdR8Or14BglwOyTHuxX3jr9ntC5Ef3ET3cuMlYc+sr9XWbG6bVA1znyOOoPnMAi//
HCon2Ss+4vrzaKoj1c0VxbwrgzPycdu29raf691EhzfPz/6po6pgY4mwXJ9ha3LA6Mjb94Bibwf3
Zx1LJrmTzBPH+DBlDrQFUC9v9iigq0U4o3lZ+Dx1/+7iKdo7mSv9tYkzw/AtFsUSam9nwx0rtVon
ECrSbrRh1nynUiuLMYVEsH27rOTdO41PEyOBupnQMsFnClCXYs+3CAQo3/djwSwMQItH36s2M5kY
IBxk811Pw3WdfDhR8KaKzHpjM2h4j0J8wQGCs+dAh8ldeTMKPix1IoQZ2am/tXPv2q9OqYogyVlK
ChCzdxpOdKdMe9cs8vxPfTfDylQNX35WlAegb9hp0AALiefmQ+M+YbgqoSiyy0cR3ckMEJMXgM50
U8nO3YZjhuFkk2pzC7o+4scvsNJlo2x0gAi9CfNh0Wxa6WoBAe1RNqsfUhMzGKu12PiZXGCYxfS7
V3bOqMhTn8vlC3AvmaWzl4gTueTjum/nvcuYpbTgdsfje0wVm1ICYdGJiqcTgPwUM1D+Rv+6ensG
IjXUyQ5I1wIn0mmAEmDneSOtlGJDfTDE5Hy41XuDzxJnt2Mj2By/btMP37iCR/0MeD29ANpeDs13
sONepJvpSZEWLJuyNd5hRe97YNVoKLbJLWFX22rREujA4dzos4O1j6AkPQe4EOf6bJ69YmTOOKge
ooC8tGoeJVeney9grWhZCKD1xMTBFbJ3vogkrz6PWQJbQU8fjDUZgaTl99fRxa8j7SlOnQwyoZil
wuzB18q+wyrlXJ9vGFXJlU3re6EPh6/yABVwHWsVowVtg0TdHGxFUBMcydWcy5YfmEdOUcrtr7X/
sj3iuUDtIvPZquuiI6yvK/AgOH8ITBlVmD3KpP6PJjFrbBPsPtkbBQUyjKra83NHtt2USR8YsJii
epZkSnYdSyZLYpkX6Mufx1D3JZRz19xaewBK4ywDJg6+ujXdc/X1ePgjv7vPTdmyM/TTP3ItcFtO
vgrPdNttgLxypvZGcXK6go0l//kOCRu2hJHf3NmFhKBMmEru53ApUbmZQnwnXTjkLSRVcNqcRKsx
3ZuXvihz89zrou+eY+dtZVlgvhzXoNQ45XBiGbpxP6UXOh3NjYINYu7bk3riH5M77iXj1GIvvcqZ
KUYJQa0hWaBNxcwRlzECmR/9x4JNQrq+B31PR9pecH74GghCNqpYt1aN8QCV2HmrbIjUPJSh8MKI
tYdBcGWltfDfXoNdvx6Z3J5MI86X/EP4PxybOe4luY9D9k6TtpbVCXNy6NCXrmJ/P1xVOQFZsvFs
fwC2A8Cdg3A5i/v/j/PKh3spPAA1T39YISMIKnxW3dns+CLbzVlk+bEE3a2+8T0wnwmr6EFcKleJ
JLV+auceFlYT1zoxj6N1qj/8iWSMF18vv1TZF7FjPq1fz9uaXQx7FCnd6za6SfhYQn/Mkr9jCMjN
4YSYL1GGGLl84qMpZ9NTunmJN6v7ZQnpTtTCVvVVWOFlbaSEe/thXNsF2zhRjbKLou/gUyhJmSUY
FCcIH/afLPh772B3eo3JiXNDAV99fkn8FowU48C0/R1zFpTpbaF8wTx93AMokuqi4jLQ+cU6DKZV
oL1Q4pnR7fcXtgxDM/uTNSJ1lAtdMcOH/KVDal/ZZ9fzu6quMeTyMM56p8FmnkYoY9nhTewC5GIz
Kt/lviExAUMIrLIVTeuW/LZD+vpiD8K8pbIOox4GkavMKC/r9pgKCvf4QCAxjIKgVZR5djOel1Bw
ncy+Qu3VkVKUP7UmQ9wOsPCZy/cMqLgxj6sUUVuJBKggvTq/APzNw1StTfeDwVFceMGKz98JXPZz
xS1L9R/tyUiwiymBSWC9+N5d5LlZzqmAMMypeDnBJ9VO5M7jbwz44ZGq4pHkyBu5GSeqJGHYwZHI
1Zj2GYiZCBRyGluh4mjgl/Sw32x26E7luftyGB/s1Tn9UNvJgzlWEVoFTtnq52AuIR7OT8xP7QNJ
W52u7WauDRfoHKaVFeSZtUtQvJr2I5Q2MFG1QhICDJ0VJG9O8vUCjxAhrhYqg0mILoNcah+FpX/8
+fm/8tYVD2IkGrfNG98DPH+Ff1vz7BwvjMXwqJM+2alKwjsigbNW7MkHkoNgThUrqPiV7NL7VfmB
uShFo2cTFJ1/PVGvE7Qjd/uDz5t3eTYrKVCC6+Q6I0YbObe1yL2OyhMDfVOxjJAth9qjw2mMZ4ND
9Pnry6jNPqrTLmStoUwYHZw2jza5NWbHCLraIWRGKACJ9cbgHXEgmGJEgpNvKwHcvNuT3wiHBTGZ
HgIi5LzhSoGhKwSJOcEvmhpDoK8FkGPEkIjNgM8Kpo7y8lMESjywXJMRNfnA+quRwALtLhzUl4u6
JhYdQjJD8r4Hw6c3hYElL2VM7Tb3Ee+1H1aSzmtopHtcjOStOEtFczY4jtmZwUbF8glkp16rhJTQ
D/1HdWEz4KfYEUp98YwnOEasLlNkHSgli19uS7l0jSQ9geikEy7hSi0mKshohDvQ0nMy3CipwEvW
VwXweOPK3AxITFozFwKhytaHKyXILkuDMIqJchBg7sAWl2hgsMNzdOBYOXajU6apWJY5k5/S/69D
NNDhZwrIJhxX43kcrJF+3vTIzQHAWGsIOYYJNhlaV3op3lItHbB2pQMQdbUadl+BIAbt9DgfNwPD
w4CLlXwR5WFKRTDNvfzv29PsDatKy1AUNdiVsBwknhdAHp+M6dyHj+M4F8+y490MEngewkW9N+wx
APd0/aH4igzdJLQyZPHdc1lVuMirMP9ULYJCqzWrmUJi6MWLRC2b20I+68y5tyZIh7ACIpux0dOs
/63/+Nt/mJEAIxvw7kqlWKkDH8xh5Y9LiEnOoWrzxbaTo6Ruq1D7pa8anfZHgKwoCkSZvaAFjG06
lilC7Yov5E3P35VvD1Gxm0k4qXIEiPyO1SVd7jv+i2wKtVZG2/vB/ELvtJQ9agc4PdZer5gLpWFT
rGjequL5DaQIZPxV4+vL07IzdLnZOzJ/dcQAt3A82D3WTrPL09opsz5X4P14tzfAFdKqr/m+x41l
leNBImvnZcdOCFYSqCQ7Jg3q31ViSoXksrkHTszJ/XCcM1sGGxSSTunygHU1wyNWKf+/JJpVheDs
+MbfegJHghYeW/aF0evyb/bG1raULVRol678TzUDw9aXGdmt1At/1JhmACuWoArhUNNbvAEwwtQy
gso82jxe/ENHY4P4YfWvXvKbGjS1tHpqhMm2aweseJje+l0up0H2yCLZ7Eb5zjwVgVFymC63cFnT
YkDIvjLvI0xfSN02VpEH0whe9ihmYuOqB8Rj1ZU2Ga0VWAjWP2YeI89WGEG7hqwkNtEGbPhpmWy3
qxnL6z3Sb9xcnHj7j10v/gVFe77/4APiY2zQsoz+/dfel3aoCYbYyNMS/+redUROQtlduAquK4VF
29KdxtiWh+OUjAj9v/+QPbcBi7WwmG7KL/CvpzsagAFMSPZ5/VoU/RZkZ2xsvsPeWOXpUMnTlWjs
F7LKrZJg2g5czljDykZGy4LfKLCQgnvu2Zzw5nGZF2EMK3jtw9MHSEzj54Atn9RHTnnggte7IPft
6u48pKQWLMDrITULDlGOsD1zjNBhrLg2fCVj8w/6HKzPZWt/P6PYvHAnCzi3TQFyOp2l4pBY0WZ8
PqHDSYjJiFwfnGGQ8BZQruCVeDJ7BMZzjgINY9Ie76XaKlzq4kqi1FpEYhx1K/XghT2ypSB4kMIm
gq79VIiU7KYptkxxTu76XvJXeIXNrh94vVlrsqk6MQ/s9wVNfKY/GifKjF6YRj0ljIenFMU1QXos
iec+iKttOiaE6nVxBvv4XPWUr2ow2kphGU7axJJrYKzk6KrEAVdUMqIrb0rmqja7e+w2YBX+Wq/A
hD1U7Q+mYtOXlzJMFtqVbO8ho6EjRB51tXp//wuOvNp7utn+YZfoUJGRRqPE+ko1GeocxuB1CZaC
LLSo3KrhX3wbxI6/wgE/u+Itly8bSx9FyhpoZPwVuF3pyhJFT9NQK30V2svPGdNKm5d3HnLLJFLX
85fuomNtvde/465l7EKnEm86vo1etQwjbpuzPUWg+HqO7RjEmjOO+pMkCEXOgoYZgPVwmUKezaXh
MDsiyA9O3UcUaf50LElrG3rnWQaGIAeEb5ASPntTJPZmVy6fuJS+5AV/nmi7hRl+DF+FAkxYsA9t
AXea+c3ITkqCpW3k0eI7sDVB4+8lOaDtaRQNFCAHFL8uyIk5XsbEN/3tMw+H467grTrROtfeuBFN
wlGqpJSl+u9aZz5ojw1EgBAbkHlSfqjl5YuuMe70Uuw4tytTPYI2SkSKzKj9ISZrSPtrW6VQuO9p
JxxOeDceRjSJ14eIE/WFgZt40Vf2eb1UhwbxroyTTTNFbZEH+qsbxeueclfOgh//7pz5VhV80C5J
0KJyEZyMMz2oGTXJefpHBw7Kd7si6r7+rGYxvdJBqU1Y6aLh29mlRjodMEpyB8SCVh1mAaK8IT+E
8iTWhc/GYZnUwJ6m64/4kLYo72b5vmyKCMm5gKTCxTejEsq1rTBCQNevUIFG3a2v4sCUBLiExuFF
0d5P+HjGAUarC83Ux3qYdDqe61psszlTIzKNF9r/djuTvjJfsMgnhlO6tDiXbjTiN1El5BqKrJr1
kRZVZnlroIG7hh3j3gxRlp3iR8DlU1cIBcJQ6Q/+KuLNID73hrMLxQLJYTaHvNToo0JSHkGsfb3a
rOZ36CVoDQ/e6iWcwqf2BAwDiPmOB2UDN8V5z/Q/LDJiWqrX257ab3S0n63Yk8GbbVtOPD8kDI7s
JDhKMfWV3ccskEAeuTPGip8hCgmdf37B4UY04PqBeLHJW68g7h7fhng8Y7rLqGt1rFgfY/Mjv4kj
S1NkzdEizvbLCXrAs9vVCDbmDENYgQEHUY/b1cKX2CpqPTNUIF97ulDsqqqkS6t4Z24hgLn75un8
WwOH0/BxChEyZKrqivam4aUAmVlyv/Rl0wslPHkgZS4q12HePlGpVxNjJAlwbfXfUyJ+F2f1a/XF
mnNv5E4jG24Q8Gd6znrGCqYHumZhUlgyPzFobdIqVjodvrNzjIIOdrExulAmj9iXYvE5McmJBFeQ
gZfyq86KabSGLQIClbaPMkSI3I+60Cn1zipv1zAb2wh7VXMLI77TEOTdpV4QDVfs9IZUU367w/Xx
/TiXl7eKiWKqQsu0c4OCf9+iMB2LdnYx8+0mixoxKExzZrfreyNoxhB+m/SODUBP2xkMewRALTNG
svLB4o1GvmMOLkbz2Jif/9CytojU24AovNYJjsvZIpPoR9oDC6KTL3DP2rF5rIZvYA73/+c2bjnt
BTvx2B4NqOUejIyX4og9Dp6XXNXf5HzRmI4IM7pCM0glin0na6EgBmhWg1B6LBqyZutRK2oA9XeI
ewoiIqd5r0QKYs6kV7T1PZn5fV4ND3NLtWUX36AmsnIEGUdDFhtRaDyJLxbcDDYPr+zfPT5Wx6Zx
z2+xpG4a0ZJGKQf1cmdFsy4WPYdPJg0gjod4iKsA9b2pxrAoeauCfwlgPxMUlDWrQ7ud89wNwyrH
yEvQ4hZuN5ojfXLKwzshFHyGg7i/1OfRbV+fGQEb/RVF7FMrYkE3sj/Emsco+577r9FQJ51mYl5R
y8QMAxToMnm2Kc2nraWoOPDcZI3TRYuvPF+3gI2ciTzZTET0+8IhqEAMD6vJjZMMgGeXTjscNsIt
mmXfCcb/J1re/IdzSVVQ1/vi7QtdFhXMG4v/DTjNzqNC7L36RjJqu304Vw65FDR74QmmkAswVxRD
rrHtF8BpWd8b6UU1RdNQ5syPemz8fy590XapqLa2ILFMUcmSp97zkslKdG2NkU/wsrVlBhFj6zuD
bHkhdvm8sMqtAFr0GL6/V5dy1h0Q4uJay9IWO1caD1qWuywiV/RNA+7P1cAN6Nglp6YkUP7OWhh/
N5JHhYPgzAk01poeDD9Qeb1nzB/mmq+2HT6jGKfzWqYVwjLSjnHbekkIJAOPVZK/a7GQcatRydkx
Pm2F9/4TiBY5mCVHb+FBT3uaEbieqEHwYmsQCzJ8x1cqH5eWKpBPRuNySxE6HNd5bn59aTIkMwLc
X74KZXFYJx5319l77DI+mhY/1RLF7cT9GtmeiTfsB7FypledQfffHNHR7+dIv82ZACd3LHPxtL3x
ouaG5SvkKnrnbj6fKUBE08MnzudzGhUL8svlbUW10i2arLlbFNiZPdhbxDajm1uJfi9leWnFB/3W
PIWAEfOGymEgqPLzWvxp1GSyYiv4Wx9mABsK5LTT1m7tOGXWpRlO7zgeSNa0thQppX1cboMlSwv9
MHC7X6QcBw5DHYhrTh8hKE4WJoQ6e2zjK4XDO5ZuLmTj2Yr08sGux6x+9d93nA196mNYWQS5lQdG
kcc2LwEc9+ocDcDRaKA+aoT5xCA5JActjSF+DP9dkBdNjKiwuJz/n7CuAOlOyPm6pleK69wWOWm6
gbucrYXFyTJGbn8nNQ2y/hU+9xHTgo4F6Irf/X6d0l00fGsK9mKFsxX7LGQCueI/YwEhELXiyIBg
X7NOl3LzKIh03u9MLCsLufkQQvvQYu5NC6404AY33bKN+HBhmlj8ZkjaAHHPRluM2KFaluVdHu4X
6mlmayACUHauLNndAKXCyy7ZbVs5T3yBpfxMleRYujH1/v7xuHL5azOzH0YazhsNVdd2Rqp5NVbT
vkJPpT9WivD3BUQnicqilG5rqnIRd1u7+xSzcnyKddTmxwlJLaKnM8S6XzF3MhWwws15Fk/9wyMx
KF/xMfusUUb6YWcbNl8/czZdzyNiGbUpQkQWuiLLYvynxTAN8GAnbY06agxdhrdFxfGEZkZf0nbg
rkacbmDskEHPKoAvlrDVmWEOWpqHFm9HZmK230evqUaqn158VccrbuX1wgWPcY5I1KBXfgtX5UOM
f9GO2zs0195YtEBAqXXNytiN3cHtWXucWVNgcZt3sAhRDVJC3hCsnXwJww4L4orLwaa4FD07Hrew
q5j/rKGMfX4E8rR+oabeHl5LvlInmZqiByOEb1xSalvRYCythyFd9X0V/hTIAXffR48TZiw0uDEy
imjPnfRjvn0rcjSa8CW1G8LPbDPBjrGrmJWjuO7Bfec8Ysb2ApWfomgNqPugBHARAYyehFOEaNx8
Q6HfunqjgKiMJqqjMYpNPUh62HazJwNub47Ny3qM1APxatRw/QDP/S0EGXQgf8Y+BYH83rI3ozDQ
J6W9LftlweTnzHa3AFiEwGTv8i3Kr1MuoYHWA6IxNrYd0q/AKHf5Hi6mff0yEdO5darq1+MUMQTv
FIQylldp1L5Ups7hdagqWkE22//XmlOGS3DdHU/+57O2XczWAceLTtlMfJf+jsmpTlXCD7lBsni7
jRgIrveru9fVuB7DDoynWNgbyIs1gwoOK8/g7CRmutZC0FJU/HCvD9vaviG3IA/w/Rz9c9csX/Vy
MWzywwt7d08bWzpx49xt3aIRAnyrzxV7iW+2W2JHLwNOXr2lCrW2tTwgpsd/OEWQ8UQxLK7A3UWU
dT+k+R+oCjOI/o4NS9wLNQI/vcbczcT7Oi6JeAaH6MZaW1dtiSH3M1+RvsSABAcISGHA5KoT2gas
yGd8gAEHXW5o5CNyMyKfD1LUZ/HItj7edpThZPrzUYtr8OThUSLTEu6eyhjkuYYQxo5kc/TrPZdX
VdyA5HviDW+0ydlHl5Fx7AT17o9yC8WlDbpT97mZkL4YvuGXNqzinQGKA4Ia/MzLegX6O+pTEyEg
WnlqDOxhg0eYWqw9anHAk3eNsVhADKYMoy2RBlgi1kPe4GwwaSqictbwg6TedMcCTiTpN3nYsjEA
+3y0t4AnaLmBNbZusD6cZtdBf4Fp0jGVIYe/J3p13LjI9KiLL1m92/LaDynTMfQ0nWpEA2ow01e2
mDRDN2RVf2p7JxE20XLe7/17LW9Irkh0o2l/5CauOBgg1eQlSa8cmfuf4a206FxrxfogyVmV75TR
XPorVma5+AKU+7MBfS1Bd3m0w/m74PiJrtY+Ksz0whnfakcocPW703HyN9othy1tc4bNv9qbVZ5U
Z7tLTTR9zDwE+TZIHiO7Neyxgap5LRXHwjHzkiis7+nOwIJF4HqzEMaXbDFpZ7TDxl7Eo3jxsghF
hFa9ypoXL6BguYycD61UECQLzQqXsbxzDWG8tMKUoyvTWIrNqMLz5/ElngpzkAG0TburTF5fgSpd
xULGUMMNtfSHJbJLmnU7zuBI+AGxxp60juexpyJh3XFkpRR2uYJ0WOoGSBHlCFj3qi/k1vqk+TFn
OoXARWYuAkDB3lzIHvS0+U2IWHLKEYn2ahuN/lNDbR+zKecCt9BqMioqTlktYZJS6U3lTz0iUH5R
StOBrmvVhScNCJbhQEMUq2B3Ux3UC9tnqHM/cUSFtaZMhOPOqfrY7tNKwMslPAL7uPojjkg+pb/f
hyARwQQ4eS6i5Cw+tXqBEqkYmHjgKB+UdXrDk4MhB47HjQVxesgpMP4I81SEgIUFUk0z6VLnpq4I
0c08FVpf7Y6hQfLrfuCgTMmQQp2gk+EFsThMRCrBqP1cr7u0jVpW40tnoHfUJczv6TvL7UxtFYo3
60PGbPUJolwENix8gi7SehADeMG3xsotlxXmbAZjnvd2fx2y15CfcXtJUOtZGYUqCi9vi0iFaVhV
SxtZshLKbfbyn1ltg5Whk5RPeEG7pcu+UjosiBHTAXr+ybb3x/F4O5g+SzPrrp2fl6IcXjSYTspt
nqGqazln8TSiqoO9Q+E8a13pFqZyr8wZeLlsoBFNViMVJueG0mWO/mRz+x/NTaRSaxO/Iw/gCEuY
cwsx2sU6Q+Ith8rrMDl+BojFyFpwWG/eGXwxtUuHkWStqFufhUsETlJMAkgbPPSimKLsPMp02cqN
RC2FmlugIXwkwLooc4X/TS1PbkpmY59iR5/Tx/3qY7YaE/jCFmMfstNGT6tQQToMS/8anRIZBr04
tJTw8o8clcdmj5HY1pkuzqwiooS3rdmVSTYG41P9qk1OH/4Q4+reh3UATWrHjWY8fdj8PTMSAd/k
ZGLugOhJVjQPFcF1WJp+mKjDaqFQFL877zsrIdqc3w/gm9UCIgBim1yfSiLk5qVEDFvMqou8lYg+
6MIrxCnYS5CWivxhdQ3M5YBvaNZVOFr+rhD4fVk9MRbnLy0w51WQ99uu1u3pGKwnHUBwHr9KwxoW
GT12bgZRgPYgQiLgXsKV2UKuT06UvR0NXWBYLeqcypsA6vjn3hb3eCpZtlN6VO6DveGNJG3+/gR2
JLsb1S8jRNkAOIxrYCw7kTlRumQ77AFnAtdic+HCyVNO9ayK1UiIC3yF+ttuKVoar0uupi24x23t
zWfVQtC7Gl/WxpMjV/aA0L+7KqN9TqyZ4LgWpwc+kT6IiTgJ5qsKHOjSSV6pxyI7QGl5JU0hKUmP
maCxqOolElPnBYcgi46u2wWdGEQ5frO1Y28oJMCnG+8IOvA258Ryv1ZnNsB93/kRd6+3YAj5g0hJ
qJo3AG3vXHQg9dYAPpQeO0IOqX86I2D2mNAB4Ve0gE4gp957bmD24No+NcK0osU9BXL3iBLWQxS0
eXm/c2QJ2WFuAyJLwqCqoQveYpcMp85DlpIeHPYZpipF9c3EfQgfT2HUCdL3ddDtGhMO3seLZwxX
HUNCY+XWMeyJMJa3evWGpM/Qfu5WZ4oAp68PSXJPFRxWQTmJ/HzK1GmcracU98KTgjZzvfy0MFPE
r1kUkGHXK8cCmi+rPsdarTXjumwRl1kdPkzfQxqLK9hZRgLtCbeYDDIKiVSEh+HQ7uw5Ou/ezgGo
JmEW6yEpyP+7w5zJVeZjMIEP2I7R1svD+uCXhVNHOKXwEpacBtIo6BEMgI8iVN0IJWkHaxeqcxhR
ut/DSx2fGJ9tqVExrjszZ2HlYtvnltY3bSYNjVFzHwFMujNJd+8RPxqgELQByFT3YeWJ8DL4dP62
f8pg8wTcLgFqixNqE3HcOtqbeiTTbrous058Vslsf2CgUbZsJgO0SLm+oHIvYPgzkjqp6ffj3899
P1RvH+CdIb4DXDsMl527+8Wvan9HgQ91int2bXwKAls0ibpbLHSmUoCdqpXsjr6OQFuNhHqghv96
pOsDgVJADPTbtW1PIrfFPS6QR8kdiIc6RsvA8Z+glNLeOsFCLNRtxjMEg7GX5kPgQQIgk2eM62Kp
2PQ8931MP+W1d4A0OhdZ1nJFPGGLKPkKRjWydnQeVTbrMYP39u3Wp1gttsH0lXGmz260nX6EeIBO
wm6QnfDo1zc0icHHiTpI8K5MURUudhEvbqKfKWkZ1P7jTztYQrrr5iAiYrKUdqfuLoIfTH5z3goJ
hJTuJB8HZ5QO4bxPfR5q34m+kWcQbcf9KCgj5TI96qOn6YlQDDKbDvnGKOvuuuZ9cWgecgz42bs9
nSmy2lI9lhgdpaZWxuBH4EQQsD0/9dOl43Ctb9Yh4l09aQ7OkYiNLno7Kfk/laYePL4o36K6tSk3
hU6QiRVn9MAYPi2SLc4iwdkCPDf0FxHsnB48JRCheqnbwsc45pojAI5OorcAg5Re0ukjexxeyoCP
iz26EnHOPBlRN3uvdDYH88PfDup0Dz9zzuh7Jt8sJ0lB1XLef3pgWMGWagPjODp/uhFDtdAmvGbH
hnxunl5OIBGIhR517NGbikpg2qqz0l2RE5TwMNaWll/7uHyiMYEdeSRn7+9EBGoMTYUZWQ1kAoCU
i7cgyTS9Zx7icqZRoUN2K/L2IMtPjJGUFyP4vxeiBiFpSPC+gcbkfwJzx/OCgCYJZndus/krAZZW
f7Rqcu2l+Gg6i13VfWRawgkTOaOR/q8te34EmllY7G3HEFeIksROUlbcLp+0dOyXatPueWuUd3b/
TokiM0/0fW3meDuEHWkGM3prWNvLLNaloYMdHzt6NG3NFU222SB6IgJyD6py2GGJx6pJZBtSbKT/
mPJrgCVVox3jOy9JGPmhFW73Pnyk4stlWnq0r2x3xTS6IQZKPfgkpJVhwgddA634vFfp2YJs1CPx
4DvyF7tmFHamf8+TFSXy5KIaFjOOL1q7YV6yIIddsi0pyEDqQHCX+uel85KhbB91qYaPsozCq4n7
h4e1ETZ0TaTTdmq+q6RrSbfB3i0E6ZC1ShiWgt5jnQhgEcmO8ca2ZaXsHwZFQSgX8PDOXYEL81hi
ukv4IkO1VfWGRDZ45O1Mp6iCcZ2R9/sckEy2Q0VfWI3207Z4C0MHnGtVz6+IiORYfepr8jDeFS28
MoXx136FVUU5NyCU8nlNGdVCxW9soZJRivWipVovfP+gtV3XHmQM3KB8TAxka+cXujQEB79GDp7O
+sJ/UMHty6pA/eKp1sdxD1jjDqb/W77BTKOQjspyHPLrN8/k+RP1pjhXzllQaSZuWe5gsEV2T0Bf
knUoB+kz1JD28oAIsOoy/spbUPrgP9sfaTF2uY2238nsmDMpPSGIqlruwD/UdxRofL1BAi6ADbjd
KTzMBW9euMyfFb2bImIGX/nuI30jHUB8sjaAqOYtttw3jbkT+BlFWD9jHUhUxaMRpOSLgzilKAFO
TVcACWeVcCOF7VqThUg/8a/sQ6qxxywqomGj7d/jLBSAxsYTz+GD1T/3Oc2/wx2AjHn83PNg9dZp
eH7WTrVkhQMcMbwMdgmMFjy0US0lU1JKnZiGqApHbvkKsPBFVU4hUqmjpMLkDUo92LJWXr9W9zyW
+3SL1Tg12fdjZBloEuD0y56rUfZPx1+pKPh+7os6XlUlMQFFhKoNmJ2MInU/PBvdQMifyR2/6qHn
m8teMoFuP72DNJl5BfKhnaMt9lCtKM4rFd5moTc4hX9CfnslG3SChEHRsA7wGlvn3DLiqRClizSD
432g8cfXcgHj066IkaXyi0tjuxKiiCiloVunNNdDBkdT6ilsSxjhT1by2SiO60gYgIcV9M83UEab
ukv5w/ibvU2cGM8EYny6avJFO9ftpgTRdAyjQdHK0QNBlV+8pE4IjQ5L6ln7dMO6UdMW+uqzHN9e
UfPgSLPFTJW4r137sHTcu1mYWWWKRilLtGk6rlYdX/7DsJhTPq+iq9iWmccPG5cmCjqPLmZ1WpF7
vcfTNktdHr03xOnWb/9MvS/PtyJOArWLbIfMj8WKAbqtPqBFiNz8c4psvCgOL1zDJumhFYwKsuCS
gdJyuRL6FHHAIk4iH4LebocCZvmGf2jI38Ri1Dt0f9Kf4XqV+tOjKXxqSmOvx1y1H8ExyjPGeNjl
K0sQqKOVG628O8whKhBLZJGFmSB5rmaYB9yvUphG48wlhT7J2hCbOrBPSpgdPeQSYm5pLIJYEO2o
E76hPO5qxVfcihc5QVHgPJByt/WinTcfU4Wuv2oaTDzbhVOt+GpFxzY5W9YX5KYz2rUnpr4Z47XK
TymFgsT/Fwp5dyyTC456FQyweaHyl88rBJX19SIDpPnIl7IWYofT1AoM7jLo++Y3xZ4h0KCjDdF0
XCqZtD8ljuug1oumgXKhf5hkrrEj5AmFf/j9L5WJR8HskVyAjAIrrQGZoQrJ/bw9T7uihFNAcoNE
XfFkOi9xxNrn0rRs1h7h5x4zYiAglDqLsI6kTKvMHvKxgnKgLPHxI8qOJdSAgyrAi1Hlk4QZcAc2
LSHEDrAXv3cu3MjRTc8Li2fAjYnkug7Yqfq4Sgmd1Nu/28QfjEcdkgX9CzIejDEkGEaoq9v7LU99
g8MRDVH/xPhG5UbcClInm8x+2/8Tw8bJmOkFURs5dSxljSOVThYYWba/fsS5BhIBNpN4HCZfcaTV
ATl7/01oxUccjaLnRSCayi7/pT71gfCZ0Cgl89lc/9PP6hg/8p/q4W6bQyeYqnM54JbhaCVWwQl5
mRmh0M/vIvBlZIg9fN8Jsqw/U1gqUyEpBt5mwNWbvZqtjqISlGL2ggxtY0aYcKN3ElahwUpMEXoU
oNj3cPcDB4VbR2sbCqsVmJ0YgHP9z4Bt1ZQ2QxEoAuTlhutlkwCOBnzFECdyBLM/NBvPRssZEZvu
2IK69Tq18Lgc+sFnpwxCQHK0D+m+rDc1H9B8CswcU/SGY/3BJ38SucTIL1nPfu4JeAjdTPxqRuHY
cBwzQ4g85SvXJwnH9roJT4y/hnsbcCQ+V3fsvg0ZLwsLsD1HepjjR/KgJTWWljEck91rBuFKdZPW
UPMs31hnolz9tQbV0803LB6AOBWdgDglaYUgpsG6KRE7UISLLplgCVIHUoe46RwBFPUatwBGFHRm
otxMB0fnwCvzAyx52tIYx4iQY6D09/12G8MikleeafzuL5RvGbmyZpzInMy2GLORtQhTFcxIFnT7
/wAIC4wAwv/aRl3kqXNkQryo3NxDcvDSE1N9kgavv+VVKZVw7OWDRYQT7GmdZea3QCYcPw+aHzBe
+042YzGxl9C/+V3+FnqvLVkJO2ePaz8jlSZ3CJ3syppIm4mApDOhhHFjsWFQ1xrh3A0qWOZxky3K
nKb9rUQZzez5mw/k/6PJgkC/R6SgnsBbZwo7NZyRkfkPRaGUGn/rg0bT21FrBCWOv4Dyq5e4hF0a
BGsG5Wc/wHLPNS7eogFFzkSH+/r/mipusyya1gS8cEKlTqphr0jMWbjduaTy+TMOGBpMG9PEcBx2
XUQAjdSSeL/skd/zfKO5L2gUv48a45mdv1HI0+FDXu7t6buUhu9cGHc+rOtTYt8It173aH+wd+xA
+wX34AmAVv5GArqKCuagtGrfMhBcF8WGHQQHzu8qxl8B0vVBIzdlKcTtok2qx6u8jeWc6MVWsm+g
UpdyUvDZc4FsvmAvlTA1sgNcznpLhEzmWzf4mmx1c5KKzNRdDsTSI9a1vhOwE1tYIkejh65PoISw
N0Zh2C3pYLwTzLlStbkzXoWN+jW4/6HFpDdT4wycVnDvNwMf/D3n/EjNqEoUsHlHVuNcJWUeUpYW
IfBzhtsZKjXHhYDmW5MYwzLCGF97qoSDPO5XU+PQeW3p83Sbt3lO2hsWmsLkHU6yFRC8+4jdeVyw
wVpaB028WL8l1oQHutmrgI4ZBMOAPH1gS0h0XirrHaKWnPqGcx9v+21kYjTE4nEFh6MMzWq9XA2c
mjlkAMCvyKa898zTOs5YzK87WwVvYEOnWo1HO/p0/xZ/Lb3pP44YmtEbBrmyJJNlZJUjeu6M5en/
jJu++uw8MsvMbYoCrV03eGSYZuobUHOlPLps/CD/8+xGNV974QpZMVrxoEiH6o0a5hQs2CpCAhYr
dYo7SB/sWhwgJPlOv3zCzmK1cqBrDgVxAd0vvNZy3MTL2rSfsBOUmS8w2i8BUYskmb89oZ0GZPLn
A2CGgzmSXthH4p5+AoG8vIhL9wN0u1rh6UGuVUJXjdU7qRGuzHbfwZvlFTDK4MDYB6MhXr9nxxhc
mmW7YgJ84TGoq7d2PTSjVGCF9G1EbGPB9mCq+Ip9KLP69AJCkQ63fCUaVftV4pQvSaVVWZ82Xr/q
ACd/8QCuYlmS2FsmVYou6jbV6+TzP46vcHf15fRUM+QRxNHoiKhRek9jxFlEgzzZsb26Qw1WmIAn
HJqaOFwv7jCBXtH1FZNqcFIJt9IzU0eMHiTqsWla/7IPRf5EKOA4MCpsX8U+DQnILAhbdwYKkhuO
AETYTbuUexKxJS6/tcZmjbK1wcydqJtMNslcRlMwfEW4p3rlcZZEAhbLLVQMR5bNjQpozXHv4mNc
GFvfvJ0wLWpSQ7nZOzHOjk8mATF5Z5IcLPONTj1IHMzVW9tQQqr+qqq5XVyB1Jcdx+LtYI28PkQn
55FYILKcTALtaSc98Y211oCjULK+UwlN2YBZV/gNSDhgdlBNA0ExImqrJVXe1HQzI0mPmTQv5TzT
WgVakKYpA/P9EV3EaOBKRd5el6pGurgAjwFqf6NrW6f9BbTZcX/cUs9+8H14tnhiuv8WweUIz/eq
7Mm6djbkyLFqF9iag8nmln+mTHoygiBxQGSnjXKWZRIcQV7owWS4rZMcGBZhkiEpKQTpOCRUWizb
ZOrDZEsDdZcDnVMmKkTx59eBmeONnRLxuLwMAWhtZUW/b/lnJL1S0bZIsSASrHKjMGpTsTpk3ECS
8wclFFCTSAEoSDJWq6yC8433bqLM2yEc8OMoJXIVZwEHXTN2nm2jd6BN+WHoViyXhXA/e1eMhY+W
0jLgHXbHEApDlEXQB37Q0ztwWD8UPYPA+Szq+SpiHFmw87v0eIM11qm6cIdkEbH+E3/iVQAzvW86
RQX/nPsaEcf8z2lqbAeESdrsKR4SqWO7cZ9K+kKTTEbVn8ZeC823JnCiPOAgFJrmPCkRSBO/J3Gs
dtZ6iJSrzHvAmk8iHfvb9oO9uSS/fBC+3g7BDrSn2mLXFmffM6gKMKmcItVSvFXYcakdHBJJRWyF
Fotw5aynbUH81EnC+N/OarFy18ljdW8mEXOjWC1XtMAFH5f0NaiTCAEsr3oSpETsYyTicSdFZtqx
3+xu6F0cRaqWSYhrN1osxBxM41GWfGptbD0XB2HnT1GRPXKXHRVc9KMq+oBF2zCPBR+k4U1jPOnh
yIGHoTisIk5TtjTiLXsEf9bAxNR9EAttb5ElaFRnUVBY74+q/sGMboyI1kM9Qlo87HWYRw55bRTz
8UAsoWgxp7Nbgo8v4FyduakKHvgwO1bx7Jx594JHMOBq5bGae+neqqE/RHCjLCHHPebFkNXCzN8Y
w9A36DOWzro0QujIODlLzuEbJipCjHZbGXTdZRmBxHYS0YTzzkebjWXkMEyCLCfmggQkHqRES2gS
dL2XQvHoynIUp0fp9LgaaPDf0FLxUwmJECqdM1MysS5F5k/p0/sk4/m5BW5tG9ExUEYZG+9wRyO7
3iYjfG0v83GOZOKG5O6orOL1EBiHcw5MTCQ7T/sSUYXnd5zIV5caR+62G+Wm0Anp2nAaS3jdUdv+
OoeFCEIYZJjczArtcQdUTbPCbES22VPu7oWQFx00ambnX0Sq2ucasSzcMbEJuavkw8TXNIN2NzeL
esgnc6iis1V8qnUvNwk1L50EuNga2NAdLKRg4OjJhMK5BQLPsiC4xw5hKDdw1R8243A3sj3Atcq7
9IfMdF9N9u8pTr6K+OGOa3a78R7mlDshYuOijOoKSENbs/aeipmfcaAhAsHhuOe6xEH3PnxwDHkg
CPJJ6gvleuBNqR9NCHpa+5JK95jpESXbqOWsgxa0CzKYektAwu2Z31OEe9OQGeRk/l2XCDaa2/xg
AlrcKZRFpwK+5Rrlgnah5uvR5XPonxmrtlcujlgbuzjZGi2VssIBYoPD8XeLoMHB/zSxrJnHxt2I
Go1qu1HjlrLaMpM0T84Kzj80+PJy+XRaWsPRf4I/dvpI6JGLH1lpT4vvOhCcLMcHBDmJZ6RA4jYh
c9sTHRdZjL3s8/QEXauarbS/EhSEHYGhSRWO6LQG8S445zLMKIc6UZnc6soewtvFISrGhfE5lvG5
uS9BIW2VvimQOo/OIlVGXRmuUAgmcYQKJq1X/MqUnZCWbZ6jnFEFFAIhIa4EWmTkrDHm2MUv22zA
5bfF4vl/Qx8tJVauUDLEwWI4rtcRhypwN36GymNn7pESTDNQ3cV5sn097Jzfv+4XhRyOFInWecTO
vHdGYj+9sJi070kgAcMkh/QX4pLY3A9fKzVJfkFROTLva15sdLbApVOlpilR6GQkWxS/TsxdQWIg
W0ANE/6vI1O8NQrYngGx9wVGW3FXDXht83vGnxQQpKvwz2c6Z8y5U44VeWgfALh6a4u7skUKmtiN
pPDSFK6VWGgY72+/06AFosrbbEMn6+kcbvYOeDbaCBZkQRrCimZz8Zlsyzc85YGMTWW8isZ8iKqr
7ozz1+tlo7e35asRug9L3mAorBrTk/HB/r53/theDBU2y8DdX4y3nEtnj6Hz/3xKgRQIy3Zvomt0
+NiUrEIkVDJOwrqCQrjQtGa3YgT4vAqzO2lAK2tiXINYPCqxrkvGX8vJeYjTSo2w/rTNuO7spShz
jHiBh/wtvF0+VkbySqA3p4Gq69G5usNGSoZsksNw/rj7IgW4ZTOv5Ra91b6DO3/zfdTEjwNbzKNc
fxmdqnSUYAmvMB4I8saQlsV8QrToY7cwty8NAomQhCKd1zHYo5ctisZXQHonuy5azwIOYbDQ3158
4h8CBH9nm5+VWi3wSKoAJG2gMx8xItHFA5ljH73RX/u/mk++aPFCS89/WMY7R0i7QxihZDmd2IHw
d5j3RxyOnigy49ZfvsWlgEhnbU+UpfPh8Rup782CQel8qmY1vokrBOwEu7arNC7Eu/nU9BM05x1D
7ujKPk2zDPCCmbU3rp+a1Mu0Ijz/iJA3RUwAo/ZQTfOjn0N9pwXr1x8xsluEMim5h9aaRugcvBlY
mUf0AkIv8BkW8SMFrOICLu00Fr0Aw/QhOtuueYNEd/fkY/bCQyIf7I0GQqpKC7tnXElU8d16T49m
ZNyDSvTHtBzUTSDhG1h9hIDK8CKc3DyjGz599HPyrhHD3aWB25kNiIU/78PVSEhG+MMsbeQ11qVJ
dNyQIWr5sx+gf7wyZtqpN1lLaEQaC9zM2ByRe7Xfp+d8GaS6No+wpWGkPm7ohx55RP7y+NbZmFCx
zEHi8rMNd5t98FQSpVfqzQHTpGCEIvgJpAdRnjLN14yH8Jgviild87VpkSKIsUnqIg2WMl+Z96Y7
dNYq12dMWAjY3Omi5KNkj8jwO6OfWg0WIYLzVa1wqAIBqntWCFDN3GqbwYzDsgtW/Ik8OqqaX1Wc
0hflZ5hmgd0CybtXvMwRPswENgvj/5UE+66/Q+Y8Nc5FES45lWJB1XEZ/oieDJp2QN9DTYmPx1Qj
w+ObNaC5Oc91HaYIPDzV+UL/jsB6Y/9VMmI1IC2cWfJzhRwyWfIVeM5Q16Kg+Nkv2KBJP+0h3qlG
yTeEac6sP1+Mo9ExTOkUra74Q0BbMrBKNu0VtoML9DnktLeiUxmRerCXFqEWJZ691OdqU522EdjB
5h2aRXA/JYeNFS+L02KCyGE93EyXYcnyS8AE+gJ2prwqYrrG7hGzqF5t6sImb9bPl86FWH4GBiJA
MjQHsasLm3xCY23nl1U3i2JdOvObpoz20XcwbbBi0RsXw0vGD8kF9+W8crPZUv1SKxuHOcWgFw7n
I6SNBHvJebLd0dSZRUBExzIGU3UL08qNpQMbZUBHz5yLwfcXqa7kKT1cocGJUyvOXWNSOHDGpR3J
wGNWsH421sEcn09Nu9fjF1rL4jXejstHQIrsB+vzeGTq5QeJodtfyEsRQtmdvN2Ezb8Akn8NOlvL
kfu6SMn5RYZk0a2IaaGTh/uUhzr4NoxWMqV2shHebgY6Q8DJSM39VdSs4ufUiC6+qwBVVgjNIXTe
Yf4Yy/LWjg6DsWVbXHI/FUhIA7VH21VPgaan9hadrVs71i09P+D2/IR3tgNlY7fp8foLkLsWudUG
rTVg6h0vusR+JTrl7BQhFdQ7M1hbAV7LBH1Ee18wqk6WufutRR5je3wuwgtk5v9uwAGFdsK6IP9C
SwxtU3v8Ut7idPtkn6Tafecm5mq0x9KShYKe0xmSehC5bJVpbPeokHtl5BdYPQraeFO6TFKazua3
q5ORUxMY85BKrPgrQOlRT81wO4viLIiJsFuXFYGscOEBXfK+HBCpr2AQtKRHNXXnSCwv9D2joeoa
BQYTDA28yMM97Yb3yfva5Ol0voJIaxyFvfmeHthzjBOGfK55ZDfuPn+84e4XvFd4pn4NsU+85Iy+
xhaSURaWjKivFig99k1vWLFtQhaArrq+YPgGWB+ZJet3Q3CmlI6wOrQCtgosqzQHV2X7AtifIV2K
5t6Gntyj1KxA19Uy71YWTIfb8X0mK8NKhoVFeFNMFn6OGKqDQT53tZzszyb9YuFNTxkyEkNTx6Bg
Pa9wDhFf7YSjKi113ZWRKvnDVihb1llzdcoT8qqP4g4WLVZt1jpJmOZtrQWvuZWxZT76zKVHs9b8
k9kH8t9qlkFiP/hIoY+Q1hteIHJoaGwx8pceCxy5J+dQ0RWfMkh4YZNU/C8g9Fbgir1TEhO/EDQV
199RtskU3I7AgsF5+xGcIvcpH3GRnRzN47IPJEKcqjNhCG9umSqkDO17SCXS99Sco96g7nVZdjyo
0t//vt5v1tOy2crkoDFjOZLlXgopFyD5Kq5VY0dzdKqgmUm4Be6Vf4iNuCZ1aocPQRp5apm/XIXK
FLyZmbtRiv4CX+VJtnnTnkK6WP2N2yHm6k/6Cspa4PL9ue8bkJjdgLWW9OMHBlKsdnkPmrl96Tzh
U7h4qsGcMESPo+6CVUWfPwxPui9yxnmirzqIrAxvI07O8n5ufmzQ7AB/eBEagJFDGw1as0sA+OFf
Dg9yRfBYR+9XmasbG4CcUjySvdQt7H+q3xIKcIsihFO5DN5ZAGDYG9IgK/HkwVQmNA5oDMfG7wpw
U30L0QenNaQdJCB0RTdftbbzUBcc/Mj2i5SFf6Hih/6zjD4iYJF7YAXT/WKnzY9FSgvuaZHF01eM
fZOsLybYk/CuEeSpQo2v7JGu4BtlAlxOO+zTpwxIsPQNgAIWaYDjitbXhluiUtOudb1DyC1cJLyP
c/j2swYCVXzUVg7nfHUuUY0/EDOWgZKCn7I0YrNH9EG97IfESFuZ+BJaSrWKZQFCl4brCMZnhWIf
Bct96caIF7+wqttzB64sybPaVKDEZRKwJxbObUHysCfzRT37hHqoPecTUh96bXgkxv16UTWUTpyF
y8WZOD100+kxf+VhJfXeUnNxwrI9Xz7P2E/CpdW9p4kgNM/Ri4beu+Cjhil6QuMlP3066XfzgjWy
eVs9HMFzCwz9LLdwH20YmJTk75TviP5Bsbrlv6+UFD1kaohpdgF/e6ZaUiNvoLnyfMIvNI3B06sD
cxYf8mJyjfUJqHgxmYyL2YrP30EQFtO9Tdn63k5E+YKIu6oCwIb6ecdPDHf2OXBFrJy27dH+nukU
BxIJJYllTMfhGWJ593rU67h2Fk+Vwa4WsPmX9jqZCzn+//IZghd4CDBP0BdxcHrxAfTFemOzhw1S
QlQh3+BX+oz1FU13ER315id4H2A6DAa9/jSHhOGFnyKt7h/MFpVS35G5OCDwOGjBOj2mwF8Fo+qp
VPrO+RWduuYcGieezazvj8bnRq/GSQiYnl2CFqW1JUEU8EqbpmNZZqkoIsPWHXlSi0Vu2LCsvP88
6ELZnVnC/spKnRRLvx2DTc/T8hMOKacQwdfZgetJCn5OQuX/0RzgeOaa0rQ6onDHueHI0jflvAXh
OV6yp+uVm3nePb/NpL3CGYriRm5v0XhRnRUgggA4M21v2hl5dg7oWcu05/UsOuac5O0hOgl5S7tY
PCPiTDC9r8E5F0wXQznQr591tkM3mD2XdPyJd1zdeB8fWQoAlL804L+v9sPRP4vVfRix15X9h/Hc
QYN6WrFVqwjSp/7N+gW75AJoZGri1XMrdAJO7Y20DqjH/sa5meVKD6o0hoykqQR6N7Qp9sozjOvG
M82r/pNDx4soPup7h/jbdzZBzlCFngKXekuTl1I9cJ+qdRdIFBO+M17egS9h3odwE28V8uwqgFTb
QrMtFl9zhqk1gkdkppxsX2d+YIrr9chJCDVwsNHGFyvnw4PQqnbpLoQm20R6RM99UsRSfYsrqOuH
5wKk8+8K/jlmabg/K8qqRWV/hILr/RKcjZO4Fg4KpAOmtF+Q9SO9cb5QagYlEwBpnlVkS1ZLG7z8
dXi66gk49mWRtn07xyij1P/qcseCnGJRd9K7q0EWYMhSvujXKi7/04L78YDrK8/bInMxuu3dtM2c
sFSlGq1carmLEYZc9umSN2+xbVAnnc/mUyV7yuDEYk5ec9Y87/ykFO56SYut3n3NzWzgB/4A6xbv
7QZIJAcwqtKKHxIGM5duz4o3PiYHJHedtce/s0nZeGSdjxjk4Jmb5wSUOkCbaJ+mi6wgv66KM6dI
lRbwAnV7o5VveNNo+8/tg6YwB8HMBAlZTS9q2lNfPX/OuEd8yRM8N87DFn9PNg0zsdNa1vP4Pk+g
eKSWRPGIRD4q+tliq3+MoDF04EBhVOdsL5MJs2ahYUUn8UEN/YA5m5h5WjwO/wjz5+jYEPllEKpn
4lX9IFGvWvcn/IuhO/m0aS3RlkPOGFgFd6yxOsQT9OJYNPsT4rTNGXatgVXcj+ab3Ls1l4smfJ5q
mqqHSB0Lztw0mguYdW7dALR/PKJa+6SMmbBkshjJB50JUTbYIkgNPdKR32GcHD/ovcIIrMuWJNVj
Fms7Dtftv6EdiwT3pMngwRUfqk1MElk4NIY3b1a7wa3EQvOBzk+WpjF3wfYBgMq18agf/HdtHdtP
eEkMV3wIIqMvHNzjR4sWQJusaTMfXuEqriptQBrAStHkm4ylJOdku1qmEtU1TV6jDrYNCBD3QtO/
S9d8L0ur1/TMAh3E2mHRg7WzvBvORpp9DvmtVzRRckBCiUnZps0LvUNKGnEbE/Ll0i6du079do+p
Qos+dAukt+zahhlRcmd+3f51il3o8rXH5erviHwJMXMvt9Q9n5Xg8WyIJupYstfT6AbdMAgnP6Jn
QF3FeobyH0f1QKWYDLPV0vTkP0NOPuoZergCcPw58MYpsHXeGWIx8JMr3C2WG3QrXoskcJCyehvp
HPQ43KkLdd9x02VNYFsuxp/lralfzUCmQAVx/uZHYztbgJxv4dLqF4x9hVjfF0A1c7Gs1HiJyOO1
xxwDCPgB3OiJFksLtv1KW8OJ+x/S1OsBPm+Omcg/UmIhq+SokEqDnpl4LNJqaGn3t2VRt4p+nMA2
aYFagagsDol58BxVhdMJINSaCb+YwnPtnrwHY/OMHJwQix9+BpCStewN3YBgydgi0kd+L8C8PFB9
SDVdMNPgMMrEsC8Styz7khZot7QYZNDDEgjP3EF/3evlXBg/zVaNldsBnmvmxPpJZmO9m4CUBLzW
cle0oXh1OrW5SGe3BNq5p8l7zAvwH4QaI/ht7KCIyb59kqfn+0EuuGWeWU9aREbvzJDqiONfYJc2
YS/nb5PucoYp1Vag6bDvEkiCIiG7+2M8pxVZkbEtxSyG3ZUtgkXwm+A+owPV+QzQiVvOKxVuK8A7
XVDqVsayOY6kqbTWW6CHr+IkBqdxik1FttBQdouaF9jcOOGPkL+UY3C3cexKg6bRi7nFnPIs2JmD
a0Js9PtaNTfVibbPkaYBxBgJ6Yvy1ay3HrWfWWM3Jctf3qdUFVQvyv5n0cAdZ5PrcdrUVUsNeusI
5Esdt3ZoSi0R2miTRpmvhyNzH9BfsJKoWWqXsal/7nbP1On40ISQQgvZOFy0E1ys7yeiNN5D33tt
J4bDdIwmYS6xPZn81EWGr9USUsmvVcBkv5YMg0iO4Q/JVI9G4nDSN5CtttNNZgB2xbhjV4p1Nzw1
zwQjil4mbro50Y8/9hqfdqnnoL1gsEjpLuXY71twHAaXKJ4jXdVDBxiHnTCoq8MYsTrMdhzXxwCZ
W0w5CAWrOMYkPVOv9cALhMYcg6hXqM/bTd8Snpw5nQh+PZ/CHjLRl5gxTpVKZFCgNHxW+MN1S1jr
nvRYrR8t9FA1oEMJfSBATAwHrH1MeCAhrrm83n3AqH+B5au8GDmSVX8jNPKfizBxLgoWFuALfqIB
RbmiIQ9oIF+yvOCsSUOne+nU9YLS3DHnbh5W2MoQn6k8qMSIC+QNLSpUBISXcg+9ms1PqE1x5UZH
xaWXf0cjcMIjU+HgQDyo2Z4og2ODYIbOHqenHovkYmfOT6onb1V7A9xYBbqC0MKYD+QJEVq2NOMW
0Iky+yWK4XljWo4M8PjABdUgK8AWg648EQo1CglqCuorDV2D0w2882XKdEJu5ouLdteQJ766d8qD
lHOtDzBAHu/3oJ+BJnyeMk5wnfGxXAZV0jnx/2s49rGD4giw16l6YJocZ9bDvtuSHTTQTiw3cDPC
WZPjvPquw8QlADu5OGcQwgdNCsY44dfzQ10PlNgHzWzC9ADxci2zQUEnlF57OSg/wIjgcUmqud9u
J795aGlOBtMAdlEdca1ZHNBWG0/v5aT4OtsS9xxrr6h1jctNYnPJr9bMoeHmRw2iX8ckLlH3suUw
o/fT8CEra3LjSjJkxuw+iPucdBfg8N5Fr4tbUj8yF3D4DjzUQ35VkUcuLPZHk9nGW8N+GYk2LYRl
GR8Nc/VarzqTOTepCPA+O4IbctSZeizehLt4D1GwNKsSANjHSmFwG0I6dc4G8ITzyKHzHt2icnYs
iIpewZAVfXs1i25tfsEX6w2AtGJbDlZb+5wIWPMfQv0zN3COb1igsUQuCTKOiJrJur637tt6TwAP
8F0GCKrii+1MkTExzOWpComrj5AwjqncTw/jCr2mn+Mr8vd0UiyrS+URCZgsMScnN19fMvhR+eCy
uHvkcYA00ULsjOYiCkks14vtucRRD3vV9nD4Q1HAm09K55S9lsH2xD2wg/rrqGr4LfL6lT5ktIkS
7sWhMdIAIj+f5/TZl8l0Yfspu5nruGUx2qWRmn7hHLjuh7hhiD3n4RO5DeXT1caLdWx/Xzpk6m5g
Zj2CiY3Epbl91l14U4wMwlm645snpJBUcy720mJhrSYRrWdeGm7kJiQzKkeBwSKx/mNvJqV9gVJn
PqA9PHagtMPHGAYrIzq9jP9u/dJHBKlIL7FfjZu5G61yAepH9Bysao8gTc136wtZ5WQP+JVV0diB
ROfeXebmcpY6GzA32D3XtbE03dfN4AoDdcxLKo7xvWETmbUj50L3fcxB4iTdMIyE33LtAymNeuzT
45grj3uuoWA+Pdw4o2VFjyl55owdxfG8owaxXup7lyNLQb17nnSwQV5d4U6eX0vJ5N2WAx7HEwQB
vO92HUcfJ5xPAjO/R69ahVlAi7L0gDxvKmyls6qiv7rZ7kS4srPh+Jyr1Qm0R+ApgOn5fx3qywbz
OK8nVh/1Jdm8LUQXkmp7XHB6gBVJXx9blLNZHT7fh6l0Wap+5N/DTjPp9iqW26DByoaglh+07P1I
1b8s797kB0EaZd+Ade37y3hpNbVPYQHNauVjkvFTUPjLsOWd4ueha/fsh+6YJLzpbCHyvz8+Opq1
kQ9ddOIsif3HNgnGaIhYhcTdZ4NGYaLbYbtNHrvWKBFpu9XvXthazSNba2RWqMLTg4pJba3UfOtz
ucT556C3Tjl5GSev7zLXoTNJR1QaVooaKmay9vMxk1FX77+2fmtRgFxRjo/rD1yFWfOE+TVBgGdx
gfq5CJVEvPgk6GJ1aKUWS0xk8fn+6GGEBqKsQu3RMNMoMKdByASyEjf5p9f8BbLp0Ec3RF3cv/Om
d8Fh0O20kT0LnRziE0veKVaNJzd9RGhHlFXo/eMlW7IM8Y0Ue3Q6tpp08TmtKAnPZJxed7hrBlZI
9BZ/VlwsHUVGa+7QxyCaMG0YFNaD0SHKbbVKspvtqPLsQscl6eb+weQt2MnUFv2nD+v4IercA2rS
5DNLdtD0p2B1FDyEjgyRKthUsatGQxh0/vLdrdpffpB+WbDJUbsaALBeMcvSmqs6H9I9o06rFIL5
chJZWf1qmBfQpc7H5spkItQRuunfHBHmp0ZQMU6GGv080vwEhnDVzZ5633CORUMkbOD8tS/cL9Yb
r7xPMwP9kgFjlSLoSNHx3xuDKowOgd5+dePWiKasROdUQ/Bau0h5k5Bth/2Mu8qbty9+akn6CtfA
4Qtg3u4cDuqvZ9RPAEQ4JeqsHUaozi+mEFz4z0PBnzzMFOhUtUbCYxJoNHZ4XcgZqIHW0CgeLHCC
6ZoLPDSzv8evANgNxmv1gLwpc+Q5V8Gj3AEH77lNsMuw2lD5gfRGqnPn0dBuL7uI7Le+Jcq6/9L9
QGvIjyqgKmK/7dZqUKZFXen9SFQc8V45njxBNL7K3Nm1ojZLG4uqoj9t5h3RC/LMsfgytpWIuFTo
Ksb44T9Onj3FsGaLy27ryhfAhGdFku49xFnNFvzNrJDjD8kFPfPmPBuwdb1clvClVTkhq2Bo3iHO
L2PFjJ4nhna/8UwYcpmzERcExrwjgAn/whVBytEM9Kc50il26B3ya5tn/P228lAAMtJa3EQvWBLo
QPRKYSlvm8JAXxaEUelzch1bxQadAbNjeTPRTdyFOSYETNPU9eYymZR9udo7zoX3nfOIM1sRiOyJ
KmAxP40bFE3zRhlh/FTUYOmAU+FCYzLg/nazImSvGXPQ9+4xpMeM1w+KLNliobNs0Xi1ELNK5Xiu
heEkpW1gxm6T7SdezVlnOd1i7En6Ve8luaLIQtFAIx2///QLLo2U3iB+4BCqYZkQv5s9fFdIOFU2
UC7wZbfDNoCTXfpO9mJgpdq38wHjEC9N8pN5js2bktqqoV0GUN8I652nSk7BI2KVee+r8ilS3QST
AwwYpb6d+xZMr98rvRhepGV2y9oYx/H0vq9tuFPTLjzF24udnLHDw4Wh4cws6ybfiyZDv51w2P0N
z4gvq2BGr213afCrF+gD5Cg3dRdZ7wPk0vaTNJ+hAErZfYNwjnAL7mCw0H/PMYzVXUXRT+9ag9lZ
tRYF6fTuyg5sHb6wcSTDtOKZ7Q8xi50F1HBMknwFNZKNN/1FfArs/lN6atQAZ9j6gWCfI33wkpdo
c5Xp8LdE4GlX0HkJUaIv4naS0Ql1/5gPQfYasp4FOqQNUmfAk+iwl37M7CNSqWAcPbjC8FbBw07o
IVB7H4coYuaTXZkZL+kv9VkQLFDbCq/s5lWDOnaioaulgI98REo69fG2ML6mHJKBiMIngb6Nop5c
dJuwbwxu6R8dPnGkgfprvylEwy+SapbycG4X5TWXsNyPDh3kDG9ojNE5YhVLo+FAj3e+f2NtZmPl
LNLZY39tS5r7vrw44XhR6r5B/5QPyIatEjw5zhBZx1pxch27QVUM8FBsF+GOEEePudzxrgHnTKNx
V2xzUwe9mCoJdh9Oye1HhzCByP0UFSerU+LQWaYxKk2KQmb2sSv3k2bL6eTXT4Oi10pA5pq5euUW
DchrXonfU5TgUpJfUcTJJ9FEVMF8eGWwhZHAdS7MWO6tOX5+E+KPZQmGZ24S3L4qQ7mvpJKdDyx+
FZir982DTiy4cGNVzRsgtet3bp2JwIbG50k+XGMIxHHf4h/9pO5OgYpetNj22Yw1F8R90NnGb+Wy
Wz010aV1G0vbsQ/S+mN1Xi9KAnJOcF1U20mrl13X3QQ20+MGCGy2Ogy4orCx5bXXzPx6gtf+w7r+
eqDuRcbYZSLGlZYv2IqzZ3YRO9+XG6zNaeftZ23keQ33lDA1hNcF5mpq+Ygm+lkQyu5p1ap24X+5
CsgUCU3px4xajLtaw7CwsxbTJ1jBwTCbm7VMBVcg6RLr7nK5am5v7qmm8l2JCh0sif4P5uGjEEYd
rIn86YtERd3Q/OvtAlIQBf+j+7phKB1P+A9faYj0kwHPeI7abvxn1gpYig+lFRz5UNV8Wt8/EJl+
Wf/cBbnTUcZ+IC+yNQkEDLfrxtq3UfiW8T4sYxxLEEyO6BdK88KOPySbaInJAa4b6D79dWKB6MAF
Qv5KI1F0eYYZniqPWGHUEwzQSZ0bEr5/qU0LJ1Q9I9GCPzbPJe75Zmla7iQOWb20KFunX5hCz4y4
6StQomh28Qo19azpfmA170P4yTUtlRzliS20NmMdcjrB4ZTRIQNjzXlpqmTP/a582msRQhSklKcq
SHwLv5jA8xvM2Yi9aYxfcO+CSsQMUSmp8JtoCMhKoQ/O5rmi/27mgfCARBt/fNwaPH0Cuv6yHlQH
fyQ9B2F939CwVSb1kIJMg6t4ul0NKht8uhjW04I7FGbC+SEFDM1LqocLY2n807EHU4zwJLqubhT8
RBrDMm68X7FJxNF3H9dQxLMslJ6LA5xIN0d57rvFTJMGzK3xRBz0BHpbO8rImfM6Y2Atn5pmGmkA
Ip/bQN/oxhLCB+XoqzIy3oF+s+22+2B9PDSSN2AWTakwc3MvtdFBGJrEK4iY3x6r5BSdHLUaSiWQ
KOXT/AiNOwsi1HPXYu0gE+BbyZcFvJqTw+B5V5M1kf7Shh8EGbRwJTPxk8hdPvquVs3qa5v90ndk
3bfb9Lm2lSGwVDIi5UJlUyHsWEcura3W2XPCbqna/Nh9CTj8n712c7HKF3SqVCnNqmI3qIU/5E8A
+wwStn8VsL2SLEt5O63zybTnnpIumBh0RtODI5qUGysq+hNjTkG0CxFc0CM/FVtw4PcPqADeGHl0
zORXOPhprADoJ9CJDjvI4NmvhYOD07sG4u3xdNtbqYQxrre0+XBBeRRnN9cTLJwB+wCmtM+ULUDB
FjToY+bM00SybvY2PEe97SmLxrYobTEOcMTz/8ZZUoYqhFvxqrZKaA1lGII7uUtgUG1QsbHj/0uf
fHHhVGACd9yaHxDfd+soSUM7LekvHmHncseoIQlQoKdEFqkuv6jlb8at464/UmdNhumz2U3y8a7H
zZv/zam7XPU7Bmaqy//X4supdjuIsG89ChrUJyWeyKsTCk5l72IKIgBXuv3FDnw8GYQCL7+1cgj2
RNlNmcEuUV2PNZOeO7txgh5oL5j1xqahS8hSrKwOcqAfuJ8gzKQyIN3MvKT6t835z0rXPOjIe/ZY
YsMVqNpLHhqqxoutZo0M0VpdayPYUVIFJxzOikeJ2EXZZWG+n4TaL/KXZCd9O9KEKU43JQc4f+HP
kkvXR+tAIdxYljepdrf5tdGZrz6NimNgkii/vyjCSwfJU5i0X5GqIG/Ct0XhfOWt1U0fs+PlpEOo
oE6NSI/Xzs8RvZOkzwc+K/ySRpgIZ3WvU1DqmDAJ5IxTTe+KLMggcCmYa33OYrMvz0b28OztzqtQ
OfelaepQpSsSANMYohTOQAewBGZj/g8JcTmnNEyGEhn2NhnYbDkzCaVuvpWxzmVWEyHT8PM3SLtK
oBDvjn7oG9Yrk5UjOtlQrtbAaKebZOPwtJDzQe79PD26usYyPOFom15b1EVz3wdN4qCdAx+aO6/S
ra5KEdOhCNpskSfn+nLX0iYamyCa1pT//wbo2wLHDQ7Sdlxqc4j0OsPgcxbsKwzA73/SigO9dd01
HxJOmOnVYQhiCPJY3TMqBxo6SPtA7Kx4hcH2AwyUaRsumIgG9amTA+VMvd46oOHyySAp+c1QsKXp
dXdSJVHegTIh2k7jya13bl6oGD5MJUUeC3EUgXqQ+i4lZtk9SlJLJk0WjU6c4P9CO74MLcwiF5FB
pM66WyHR70KdfId2ZYsSXFOfh4p8WtkyKcaROgQ+5vE9iy9BVtlAAmb11wDe40E4i1rkbsJJ9i4a
0kB5dSUueeY8IMQVSjA9CRuxLzjtCe3YukHZaB8pgKhvwGvx06tTMJGuibIjNpeY8ifSWH34pWPb
MPyHbChrb+/bXxGqq47HorN+St8eLA1njSq2qgXX5355x4zhj8H1s1HYrHXR5m25zddc+caxrPVA
0ASry6nquSyDqZsEDlf42vJcJPhmQH+fjhc5eyLmCqKFuyf0pIQfop1bEce7iGlWxyc/yNnBwcH1
h+b7rWzbHJkTha/HKmyJKt5WJKNxiq0iwkuJvlMT1dcnuGJCKbXPl9aHZ74duGLKJDFBM7hEEvr8
xl9U3Lfd/W8XcaZEckThw1ANW8CmsB4wJ9WqYS4x7X5XF4DtgkBBHhPppOa37J8n5OB99XPQ3wM+
eRSsQQAenMvZ1q9sEEWHmNLgDRj3H4uTzMf3jSGdzIR8S8/whGX5qKTLh64/RWBs1KHPMuVGwV1D
LUSYsBqCaMka+GnM0UiC418EhIpZhSGiBToobWALTq5+mX8TQchOYaEhaLoM9cCa4tqEZEw31shM
rbs+iu0/a/QU+R8Z66BOW9vPDnpHU+xDuCRdz8JlMZ33UCcfA2dd7gFQxH7iYfBa4acMaSalGgRU
p2VrbxouK8VppY3gqgRNogA6dXDnZwPRMtYqtkmq3MpyB1LsqljAmAs0xGEjOKxIDIqK7zD9AV33
3I+4l8dg0XdLWBH9oJpsi3NFYfp6zGK7T/nDzqtSnxr7TZeQ6DMMPXt+JtNElRNk+SkaW6naLvJ7
CcZUelQ5Vh3eTBjz/i+/zZF0mKD3HxuUusbPK3NLLrOiPPcPlkzEG4sAxr5lgtNdd3dQ6TbtNi0e
hWtBQEBAz1FpGjBNcY+1Y6Zxuxd2usU7+Ex81+5ftot6S0twJsWmktaMg3sgDoHYZWgkXgQI7OvW
Ctt7LY4DSl/1oCre2yUBTDb6GpqSz9mf1tbtXIv5BnBxGwzvujpc2LOE+vp53nJ1zPE7sPiw0xhJ
Hiw9fvS8Vu53IgMHgD5QadKIkCyWlb6gYAIGlC5NQ5SREx4qVL6ontPX1V5zGzF3plRYvNtKi2Ks
sDyjQc8tq0CitKl2sD2FuLj8QcuYGIWbFKFJZzoi2Sa+GBGQlDl+6o0Ji+9cnuuiih9FZURRCMLn
m7ShJwIpzv9JRAzI5dJoiGd3BYuHvr4VLv4Dw7KNu4tXuxGgcaS2lJevtCKqcCqOlm369pH9VhCm
V6O2YZVXvJC8tWfunY4J6l2GXt4fAXJ/RTpRGBJcs77WGBG00b5TMj5gt725SapIdmI3E6BlWwak
ePQfJ5cxLFIv4L8An/YdDWc+vdQJ+Fkr+U8F8RSQ17tLy2G16TLQEsOmxWXvHFYm5wsNS9Mxkz+a
HGhdSThB8I8/zllBOepVNxB9yWvxkp4RYgBOgDP+gIfwnAYANoOo7bhZBIhCZl/0gZt683ycdjHs
opL1U1FaG1auEbqeDK7kniWK8iHSt3GyWl6VqyF74Af9E4A5ihJGTCSHoP0o1ga2/o3BQsdN3WJA
UtdH3SYOHGCJVk3GEDeh1xK2NZ5JMhl+krZxKq9AKS3dxRjn+N87U2k9Oqzw1p3Wz+M4huzARo/N
BVArTFcy9BB/iCNkeudhYftVEv3zmQIdESopQOFF5pwxZ7amHCF35irQGDgy5c8llht4p2rYXN19
wziuycW8FYXhcBvPd/RFYK132RI1a+mX1CwX/ChDBBd2IuJatPpkZVLMgThfH2w85yTfND4GPSVz
xXKen+QsAl1U/gTAvW84/FAChmdzNvNfuYZWjSCWtG+UZCjib83tI2B4B3WQAzVeXs3daFDJIyGn
IhhN2tMXtfShuFQh3PbjJ+94VMxwbXDZ9kwqfd+Je5qpWJtvFxoUU4Gl0GTV6wq/Msbyz8XRtUJR
92pS82UwLYDg03Q05cBAbQLFoccYMAHHhYIBLR5GzoUNRzusxw2XhTEZWYZaeEkszlZja19oTLxv
svM9uim+POEssdOmA0xSj/Li58+xiC/wqqYKgJUvbQcaiNZ8Vv5MmRqwxS9IL/XGdmD7KPg32JMA
krPyTVSu/HXV40aMBxC+y+P8/iTbaLRkCiFz+PvubkSny3IZHw/ewuZbUKE9KezpRLMbPZosdgc4
Ork7sJpRGU1qOI2SFnoYPj+w8cCtxtIUewTEkkGtlBxgKWhihZScF0Rx6dLiAOv6SS/AtRwZUQWW
eKUIl7hcSgmw2kaIVt7EFxJ2+Sx6Fv5M5RlV+mra0vc1xWZQnJwGbKjsz93P4aiNFy+ftv2QkB0Z
9/F/Wf4vyR4K9B9pmQYXSpBReuIxz9hURAPnORB/4ZL4IKHMg5FLTFlfpHeHbvTUVsNcRcRFsIjb
rQgIVFWtEWXu79NbRpZvc92yzWsJuPiMdL2b67Lp2a0SdlFY4vF6O/K+I5RqI85xwwoxCvb/FSvr
Zy9fgUXTDkcaJKwZ8g8M1ryKIHDd5bd+9yinONC2DV+E4cMvOyUgNeR6BOcqeep7yBFor33/8pLk
+wwm7wjJj3uuPZTm27NV3cOZo+aK9rnd8weco872H/6sZZ/TD+G1Oxb4v0J2QVaQcsty6D8doB0r
JJX+S68vSZ/qL1ICaWKDW65qaSN9ZgAaz7rLL9unMZ8YohLUGjL4g90wdMud7xrJ6iv0mRydY1wl
ihLl6tjfId1t3ureD78IRxapjb0Qjlw+rcWkb9d+JcWlHjkbv/RYDuOoJaKuRMF6j5cUZei0300y
ARnnU6GGvE9impVujd7nZL/v5CSEUy4HmcLDprAUzG+cJiwEAiP0vuqfDp4G7d1CqG2LbKaAqrHp
nZg98fogXN1aeH0EcCHjruDPxECCunwqsrxhKwKyYw3rfIp5ONgooYbMofFG35O3GC22qZkH2gCS
bz0oXRCCrwrWYJKHJsYXdSDplGaidJtnbVcop3M4xiumYAUBTCro66ptu8DVAXbCPGwFcBOvyixJ
bTomgsUNNg7uECur+EJnXomyHCjzJwMYCj0wARhcYmf1knpvdUgU/FqQwKp7B+kzajpTmiHvR37M
RitGtQZu14FbMJpU9cT5po1dLtiZyKSPvvK1Guf+xmpJkkHax6T4+Eo8JMkaN5RQ2AS6hUwyCVES
4gs4+kLowWfnFkmbirWfVjiJ4DN9nu6ydIhaRY/BgIYLf7Va+cfqix1flU997nPqn3Yi2ty/txuH
ReWNTgR5hURjLKqySAiNWm8+9p+I9jXYy3yqzTp9IVIHIabiUBQ6G2SD6XU56Gtk8jbYBMtsHFyP
yNiMRRLJkXBRtRvuO+RwWf3r4tL2A4X+VBh80A7S7t8mosa3iCi4rPb/Q6iZro3qXqjx7QM7+Cio
JgGGouxNeaHzURvmvP12fFnMJdeDozm3PPaBYu4DPC7uis+DzJ29frwUzMVsXVwhRpCLf2ER1jwA
bMD9+3g3z+IoJyHliSID61nBHJZwVrCX38sN/wKTcIOKWfnPFD1ylt1zgGYM3YCOLjMsko84bWu1
R/79320ZpoCEVM89jxz45JyeNoRUmExooGGRtDRcM1vJ874FNB2kMynLF6cUay/d0B13Q1pBC7+y
/gaL2bioTvAPUqx0rZ/uJWqdGDoPjTl5zcz0ZQk45zk2SAPe0OHcZRJVLBueyKXdKWVBoQ/zk54/
dm59InwAx6NVmD7iz5XURipjlvys0yMkPpaU0Hig6m61IPKSEpPFa5VhhPaQJAwddAIgA7Kro5R+
l6+bgVm2cfLkEr9dqhh/x16GK3EcvziZUyJxO4FeX1s1tAckNooGxd/XMnK545fY7l/NyneARN7K
32zZznd2Ij8Wha1/Pv/By9UEWNjUQVdSIGnSYf3uVP75NV1dFK8JaLIDdUMY6TmfaBOIlVhSZMAb
MwUU4+LLdeQKE8xqSayEP2k5O2UBdNAiZXKr2vd9o8DZyy9/UX1zcB3RXYOmJbFVxudRXyW4o2yO
oMso4hNKj7GD3m6OPGLjNswRI9DGpe1EN5zSauwli6B6FJi9Mc1Kma5zmuzeo5Uv7j1Dlv/a5p9t
kObdMWPMaDRnvnnzg5m8C2Flzisg8YNnKfKtYnu0XXujNTtfER+acWC+7/YZ7rWfwI94HBNGCH5L
aqFgC0aQDIdD0ZBSFb1v7sbdXYPJUHwNczzgHd4KBbC7NOlN49++AtR8WDS6UcXIpFqCgIzMBTnR
2LwapDuUdLGysrYRzAXiPXYW4PtCSLo1gVZTueJrH4tOfTt0E7l9e6tKpbeijPDwhHZJ244YriT6
OfFQOVgcj88LvX1S8f4TSYBi7VZSWPIbtpaGGrDoKk3NwbD4wnMUNTNKvC34aywtwLHMz8I9lbuy
XEUoPZu7julS3+iK7vSS2XakLHkvP5DtqRVo6b6bm6spT/I9G+kOKMIJQ0DkhhlEZ3kxRpLYBR6B
x4VCrT1RWh7h0jF7HBQU+2SFPrYQybNxZpWRG+HmIeC4iydTNdvqS4Kc4c3DKaNcI+6BXP0/WVzQ
1x6ryDNsd9oYdz1WjLZdMEX9Ga/Yz6QQ4mtFR1rQlG7nza79jCpo+kJfLlF46GeQ/4s03xWn0Hl9
+U3LReyEb3xlVsaPKhmA/x3MI/vBMHRkb7koIWcIsOKULdF+qTk/P09wcZS+WIEMspyTOzUTDGVY
6oxE6vF2XLuyBgQiwk+R1CBLKs1l7lckNoO+/yV9ZzzHJhZVBTZ1LZqUTBAn99jPyAyBVAjL3pZh
7s+SFJFTfuMGESH/H0iD/LSFbamt1vZjRLv+dQ2ZH1wVqDua2qVizWnVIgyvwSgUNZx+lmdIp0Ty
4eQmUdak+iNW4cwoaQFcGRDfGVpJPceuY7aXYO+opSbfW+jP2hNzVyxfcxMQO4n6254tE43L8E68
hpOJu5tEsl2Sz7hAeIvFni89toukGS4Anw0MTWhWPJSvlu5yR//yaGuZWHhdPZ2pREAfZT7X0MH2
jGxyttW/0KwftyYTC4ErUqtIjttjo+OKREDorOhV11Nm0v3IhCWcqCxbvulsuZVBKzvyDbjK4sVU
Lv4O2fOAXTvLQ9BHFPC/yHuerYIAfrai2e+HD9yz8k5cjnRfoF4Rk/nreA07uUJfww6huByj8XwD
LfF01lPIBx/mpmCmUW+QLUH0hutAB7V0673lfKsOlXkN7yOI5Q16fZDNt2ERQfpVJHgKacRKBfMC
xPxj6NLVUhrkt4XJ8ZxRfQG7BVlnGeW9LPVuay2X+ITB57bp5Ukizk3omLEMMKnNLDUFeh1Tumh3
5XoUp9CGIvhG/pZ6vCWQrMqhyADXB/6XIhAcfJLphI0kSb83hxvm1f38Mqhb50Os8Q3fAIArjZXU
h9PVou0cSMt/IsmNcmv5htUoWRtZ1ZPbaBnyu7r7Siz0O8GGXZY4gjREhQhKFV68y5WGaD5HRKjF
5USMTIGQCqbdUXhF89PcVvRKNBcelqIAF6TFwEnHtLeQmDoQrboce5iUCnGm6LhAfix7cN5/y3ab
6EwKLrGJOgu9Cwlg8easj0hQdYXKZvrHAtv6VfsZWJzJJZthITSi864jqTCG9vt0Cvy8fvotZEtm
f1Y8uzK85NFtkqVl3FBYdZrG4Pqg/q4La02xm54hobUJH/AAmxk3jzfcr+Ukir79jlRrsPX1vOuW
xYoH+DLutYEriEpFrXFr7W0uYPe5uBW94mdtnmb553omv0aWsEX7eCO4ycCC21ZBgEo0TuVU4Z7p
mRTARnMgpsCuRhaXyXxXxVkGrW7gbdCQf+1dw/umCZvu+nHWLf8pWisRzaLudu2n6W46RZCP4I8z
zPpupyacYQLPTlBlD/uwjFiOaKoSxqfGcPhUL7eqdxv38qy+3gT0O/+19RkzhYg8MjILi45vxbwd
94rDMmD5YxpvC9uaSLH5QMuUSOuqGudjb9JcJ+RJpiBUBZt9Nv4MsQPdOAM2VElDAtdNnjax477w
DnZo6726nqGYJq5j/gKzkJ+yEf4qHO0Iyc6FWISD4gKTc8u3cflHtQPBG2okhh/5HHyubiAx3fXw
RiTXLRjEb71pZzAar1NLI7CqeHPQf8gfS83CzYGagzWu7Bvkfd8SzLydFUVFYj3aeGzNyE/KfdIP
qLIB7KzUkyoJ9aB6fTEu3a9CyL4YwCLNJOybW6RwHJ9gI8mgcRYbKZon8wBSLrlB8UGOVMRMZg3Q
KahLDQEGdPpsGxRLB5fPlKa2KHtR2Os0Kzs3bOr88VL6OISFcLUliWYULr8MnDqIr5Yr/NzwYwt9
a8mB8FMZ4ZJfkFt/lv4s7MSbBDf2hgtJtAgR9Ke3ifwJWPjp9bOHywbi+nBdlKiVV4q2TfIcL8bT
pnzNfc1dcYJHOMkEnHO+WqtkJFO6pCx7KRRH28uMMdSPataJ3JW2qz3Cs4KE21PKW1mH5MUoDkmQ
jbRxidrg/mUdNZT0W7jSGKMzWA+QGfIxojHAxxClz6yJwkVd3zIwESKNLsEn8KV2UWv9IeAwXl+W
SbCwPryylhy3N6qsa7SatTpqngFRG/RzaiqU0zCseEgRKUoesYnAuImwsrMhIb4GvrSM3s/DY3fo
vqN0W37VTedKz842O52sZm/vVTgQ9u9wHNPoCvzH3fem0rY7C5p+eqrDIBVOgMpZtrsOt4Sqsonx
pqHQ0AJUiJ0VmS/fyL7x9HWUBC8q8/1R1nAbnkR7WvkF8CBZu4/XWnpkSbeum90FcfhfecA6gBC7
u8zfzpu+TXvp4MCN28jurtgFaQA7ALEVjVb3JnWDavUlVkxzfsiKagWWnTkY61W13uxwPQJUwQkF
OgyhYHa4lGEzpk5OF5VMGyljXwc64aIJTCtCYC7lTwmC3dWfIi3XStGL6I/dnAw8qaPe/SvliI31
e0tVBrpF2smxf+0gozPBsUoHsmwtyVusAoOrXAfy2JZ87QcnQiNrlG2UFJxO9ybnz92WuhrNWv4Y
E8ExB/XnGKft8sWFZuYL+rkLYX19qS4BCiXKxPw501cqf/XeLm3VuRRhVk4uP+7jUGf2mI2ISqjH
bt+OYX7vy++1nS1OhOvvjYZk5NRFVb+Rf5SStJf0pUKzBlVbYYwrNZOdWQ8sP4MvBPEiK+A0YTzR
yVBT0ea4xybB/cDM+yfliFCMgzbSRG9SC5nK5oGpk8M7An7DJ8kpBSNM5AxNF96SZYkIbYVHYeQt
w+FKK02i57bisgDe5OHp1ePQOTr+N3OOACwnL6Bm7g0NBN+8yU/aLv7I/paVf1OQ8JjKSmWvprmn
MsN5TO6ifg+ieni/p1Npu5cXiI9hU2GwwCla7B9fT7m4D09U2BCRq3lv6W1qTvRYdmZQdfzeQfBS
Cw9VhTmMGyJ6Dnxes2xGi2PdwX/YNMYQpKTKsb/gmpIa91p1qeb4Nkv98uADj1fAQnTyUwyawhB8
bHoLKO0B4E1tMeVzCeENMqnoX4c0drEZLxz3yREcTlmM6TbDoa6CwWTsYZTBY2UPSNuceTm4P/Mk
lVwqoyUlLypWM6gaGR9x81YDxMU7MCxxiq4RpXCQ9TYbfXWI1ae9glBGNwfmSfSfRSdoSDRGwNcg
+iy59CjqlgxJ1xJgF1wl5PFT0tS3oZKBIU7+hkYOgNdwR6vYBtJpaYdOOIets4v0eUXHBbNytU96
O902l5nWJDkpeQdEVRmNFa9U3m5FQhuYTDgrOxBID8dtmr6raLz8PVRAxMRfnVUj8w2bbOSieZAe
iOlL2nGIKipnTUoUR96223W/3HgB7GenInY2PjPo2S7ZjYxyb/vv+O1gF1X/el3ffZxPvA4WJ9Pe
tMHcb+xThlZGQtfz4ZEi/agnXdHLdQRRNoY6OiAm64E1cG7VFxL4vO3v60SnTDe0ZvXPcN6PS0ej
ZyHNFck/h0zMvl0XldHGa4rGb2IVMm5J6EM4NeOXfU1J8dn0UX8AAF9Wq5h0H0uaeBz0393ftbFU
3N9MRp4uscCrm4NvCcOzYjCeh97A7Q1zEYD2jR5g3aNEWp5iLoVmKshbvTM783p78L5Qs08MfXfJ
dBHEJmj2L5+xeY9mLvFipEja3D95/HoqsG+nUpnx7ZUpMRmpLTjHiTzVeXm2bp0xmgbUSFDLjDcq
U1mZjIx7fkk3SxfiN2ns5ISsESUnOS46bEzpnar5pvjT+zviN7/rRP+PBOoldUHMq/FrYVqU/5dL
D+ifO73Jm0fJJvNFtbIlFD1QLZKvxDjS/9HSltdKklNSGf0QmevRLrWiPW8lqievF/TZSiTcgDPi
9ibzBCDep4RXAj9AeCGRJNmvbPKMV/JvVfx2K/zuCOUR3wFvMcv46s8bk28X2+ldVBkXnuU+qwaM
WyBEi1V+sfaIgfsqVsbnc6JgegUuMkLUI96XB5/qVLaZDchKtbpfPgkdXjcO+e8LWZLjOT68LSyu
z3OqwdhIwXH7euWA30GTUimZs+TDnYgpshfxRHsly0wGa5IhV8ll7PomiJS5DEJ7gm/e6XpR/jgi
IAIejHdBfmSm0/e1+WQNXW6JAHTrezeYcq4bhqAwZcvy7mz8t78aw/WMmBHilhjEISP/2AvZ+/yv
ZraC1T9fobAMKnAitgrTfeQ7lxd+dHmi8fxCnjisUUO0jgxFe4ucnoB5Hc8vNUppbSvnhKkYzr44
xdeaZEDmthkzbabKkGB33SvR/o6Awba5L7jTI1GQh9PzeWDN/wD4nbB1TLgWHNzEec4bCxUY8LLJ
2BPiHtoyKGesHZbGx/QeZwz4pRaHOf+B8ElpLrHjWtRt6OuJodsDBlVZUWzbPrvYFDGPXqQOirzL
lUA5GGkc+FfnCXv9zufpVA6LX4qz2blKzfebNaJOOQXZ9BFkpXjfa4lSDSSXTxwYoGWaLDMh6AGj
863lqGT8CsU5GWjZaLIe/kVNZKizPAOH0tzFOwvsQAW7lvJY4uie5eKZ1z7Wt6G+DwJqOA2lRJn4
EKg0nln8A4HmsKpjcUKbFbDuaHND4Vvs/TjB+6P20nAQOtH2IgLS6M+kI+gckz5HbcSZ49jynLLA
vOJ4s4gY67Y5Q35DSSfgs3Ls83WxxfE7FNlK6kClbQ/jcqILPzR02/+li5MFD+SmOc3H7o6YkIgG
sf25beSI/YgF+J2Vl0xb0TwbtX/k/d1ZhErnW2qQ/g3GuDMvtcUp00G3QF93JteeyASt++68qu+4
N7SnpJ2Ohsp3vxor8lS5ZFdto+ko+sbtoAsRqm6NU1/crQpFL12VH+AQTD4Khn5S3PsszTZ5Zdpe
m59ZjjOOjJRrEkDX6V+jeg7JW8TXMoR2uGWStMxgJgTeFu0XqsFynwR026KsiT1/3KnMNGvHZFvn
PCPMHTa8oUGGEGg1MqYad97/KjXRGEcpXqJc5gmiEVYXsbO3Jla4zeaNnohJfnSS0SXJQklCfsp4
5+ZcGGBzjfPsk5m2sTsxxvtOnvgqXcJEn6QE0yeSj1fsF7UeKwZjZaf2gl/KRneWxXqieHDv71RW
MRzuqT0C5URK6mXCggrhDYq/4J0gzgGGIRk0/30lye9MMJx7vwGUdOfK4/77+gEYQkNKu/XmJHaZ
SuBzTF34uvnG8QG3pYBEgsFYQT8HL+KY0hLSOaaNl0/i9KKSPC20PQBsRSkp1WC1y5SrY0+0Xxy/
/E3TvOmh/xItCci0cDktdwWDpx9ZnbLgsGyVXFOIWMgkrosLNU555tDT37VLCc99FzBMLZGujl6a
Z2rBsEkCV08LkHnKj8gIxR0fdV6RUr4sWbfjAHChIRzD0EFoeYPLg0MvGYOIoMiKSoY4vD1Uxglj
sAQP680vmy59306K+zUy1dxubQwx6G6QjGGPt+hi781R70RnRmLxD12rkDYzxlXkoLhv/S8cPc7r
UD/zJNzl7xNAditf4TvzAq/CzwcgXYe1Ct+gug4QT/yprJUHRC/mQkFGjk33+dJBy7FGAkj4fPAQ
LjKP1ItqAcHCKGBUKCB1x105lmYbIuXQWEZmtTOBeJ8vAaTiPMZIuNeYFq4820S5gA0jPDUgP9lE
UPDL4Xz442TLawWvRuXta9mj6+tXZhlXasBsZADqOIERHn5aCJrtikqZhbRsf9oeUgACrC5SQClM
3fAiVtWsFA4hKayktrKp+jrvrKwZixp2Lzn8ciMpDSD3AFvPsn0Wl4Z2Mq50qXRzPhm82nNPzG7E
KLF2OvRfECYZFzitLnb5f4l+SQWTA6Juvu7ZQesBVDRFMe3twjxlgIx/XBRTA7PftUAnW5b+eCrW
s2XRSfiVdFy93IcKlQ6JclCXgLVtu/MHM3TnARUiVo9fDXvmyAI6XBRdZBc5Xk+PKJGuAwGg7zx2
i2wbsM+inrm+A2D0agUnpwWgHRIHvppXjKTEosvzgUvWdjPxBAElsYxXmFSRxoWyxuMxKocbWcrU
PiKT8l15fhRqYbATEDeRP9TfnEkUgVTnUaoCogGAVUL6aHl9HVhP5ALAATHSWl22q49aB4fJRT7G
QVlRVVbHWK1QhD4sHGONf/K5W6tXlgrrQf2jpG8UYsginqzUOXIGVWB47u/NjrSO2WPGqHPxT44I
/eM1hNb9OZk7PWn7mKo3j5lVn/v2ZO/qPW4zMUzWLpHpAwzLHZca/hn3x6ibHLTeoQJ+vEfxfZQX
5VI/REM6azX0KRRp+vHtWQ1JlwJ0zyNE83dAjo4OuTH4LODGPStkqT7F4orldaShwy7+qPdB037+
CY1cDVJZNejcCkpvdxQAd74iuvnbm7AAjW05urFXCgcr+GzzxWYs2aqyTWGhmTv1MRwsC9akYqAf
571vTD6ImrDUjKbXk2RmyJms4iOrl/e0lxJNS4igB/FrHq1nSELOE9Y37DaSF75tuiNel0Yq9pn6
LNwf8oRutAqFoFUKQLj8I0+Un991AoubiiPEBuQbLXQopTo2vJAJ/KpOjRHdTCilA/2H6tZi+KcZ
DpOOZnfFrJaQYVk+brsIzD7hnDf2oLXsl5pvU2Z7g683YGCHE2BBbRHwoI3UiaZ3cRnk83IeRLTD
Poh4R8UzsFmWqMVn3Ik9XkPXzNPzkVIquLN0bQx13EzJfHm7a/+VFlpCC8jz8PwvfOYM4/Je1bL/
mWxUQzESgbUl5RB1BR5UbeKwm4TYo1eo+8IoaGjLX3QgBGStVTRAx+z3hSuuWrGDC8/X1dZwXFaG
n/1LtKfSSxXfFuaTcZmtciya4oTTS6PEW0pVla0G3ZQX8FoKpbElbFtkGdtPUts3pnj7v/r+Pma6
iYEfdr+bFEu4lCD5ZK0UZY53aMY1J7gVrJB3aV+ljzdGtLp2mWZ3YWJldVycghKJcHL3M6IKG4Yk
SzihCP7xG5l2yGmppE131oyWCfxoFsw0VmDe0DJatIuPaRhgen+OLRVZf+chOzVJe1AEkfnnBycV
5E/HC3ygQYxq6mJCEacx+GRUY3xerwYEUE98yizLi/tmmCJXl/sMp/abOWkcqBrr3jq3UQAM+BxG
UuX1SJc1R6uJ0g74lOjbJ60Ijsg93+moAwOgN9AecpIvBR2ksow1i7a5D7bn1M0BWEjmiHvL8H7U
LZMxaHYtb6ZETBDukdhf8zdDF08qMqS/ezVfEcvpZ0rcZycBT4ZoPA6LDqEFOeeKE1S11ZsHqSM7
KziAHSO+gA3S/H7IJQd7g3T/IJz7tO5nu+MG6Gaq4fwUiebeCIC4VDEqQ+nDBMDPL/RUge9Vqqa8
RBH0UVHsUH0WVCw+0NiW0bEZGc5yIunGMTcK/UznoB2h9nbSHyxbs+Zn1G6kmcgmAs2TP10AfQs8
5+65TjO3ETmwNLE8yo1vxYV8FsWgOJFKH8rpiYHvQsPnTGAf42kCXpl0hc88iUZlpCRqQ5cYF2or
wyoVCzxt46PfBHC2luaajbUSbYrJpwaSH6YIt8Xx74nHue6ZF2/u+Wwb60uz5T3F96JzX/raWRvb
HB7EziNKT/Uqnr2XjrzkI+j7WUMC7q7ZatbtC/bB0C3YL+WgdoE1WUx3sszrr6Ls9DzA/V8Ftd7Y
4tEwYK9yjUSarbl1jOx7mV/pu2J8ngK4eaLpah/9wHtYEblf71G4yGqoCkGm+3xG5bhpJA9E6KVz
z2xFj1Aeiu8DPP+/jicnB9bC1NnEKqQNiSUcgY4z9UDdzPVg6KjZvHVetm08P8N4HkN7hPQuGTTz
/FfrTiAt+dREmvew3Oednf5E0KenpMKUoKn9tZ281r9gQW584c0Q/42gSqvrYkGBdI5ptyz7clnJ
vbZ3gtjC/SUvY/N/DpF6ld0RTS13VN8M1el0rZyFxk1Nrl/5D9cYA0lUhrJjhd+yQUdL8kkXJJ3J
BFxjSFkDkcWXMIr9tEkKgUBGtDLiSLzm/0jPJ05ufFv5VX+OVijrw1mYaGulQU4EFd1JbeU94GL3
7hVoQD75rUcEPGFtkBHqy3TnPl1UjhRkbEbsolxmabr02WIkXrGEdfhYLomSguQd0SiBKp3HjiBT
QVzxDCyMsV/khevYNbv03oNC+x2ode9Zxg353LHTXi4fJqKZNJvQAZueWVm8cAomySUq/Wu8ZUUL
WZcrcNR2GzCTakHxrCKiWol+n+j3Xvrv6iyluvbMQGwQaDGoPJhVhzX2tLntkcq3CbNyOU05W4ZG
yNja+rggNxwJNTQ0c+7zXj+0wx00mFkFO3FgV4OVcjjsb4zjNU6lke/zdWbpVOtX/CJ449Yh2pzH
g2hiPVmyqbFv1bcvNClKH7lAwE9CANNJM3lqWxAajtn7Hj4T1UmXj5ZfmcRheCcPkZVliz11kEAc
smKh8djC6BeCK9f9ZyvnO+uJBPpFohgoxPhgyKl9nQeotbroVkcczGIAmUBEsOQFjVRf8yHHCv2J
As9+wvBUVeF+cGaslnhAzI6j4DKRKaJbyRzOs1oTr2JsTSAmoFvZ9KWTOmdix9PaSbQNL0Mpu0FT
EpeLLj4NtaJHiV5JlRswE4xp+B2lCJX3ZpeejccUoIiJJ+voPix7y9TnTi92QNg7Xri2U9yAW6VV
jZaFG3c6OQdLfPHJJTqrKBQZYzBBqZIbcNyvNeYLmxRg5IN4NXP04AGwJTajN6PWMorx1ECoO0/T
B6Q9YP4QirepRus8fcuBU2YSFTXxWgZ/94jSox2ZrTfjVzYWC7um0u4IbCfKnNu5LwRrnXXstHaX
CfCAPPOSUIuZzQJ5dkJmeFMgP3Gi8EVmPDHxVda1WGDvmhGlL9z3ooQAdg+4y7cFea3RhvME9rL8
PetKCAxDp7z0eQp/OC+ydrGTF9IoO0fj3EQiRwbP3ouKZIAFSDEOZgQMmEWtkoV+3xT/NDOjfdED
QgdX595m4v9G3MmYlwiUX6xARGH+S66l5S8zTQd+zCPkJhLWAcFf2GVCxsDZcctvO9HGHFPlBsPT
/7EVIFLjtxLLi0oLlA8TCt7e9Ddclw8biHkHQRMR2ByjieEaYtbAJ4lDMZivzHViBiEQdMTvW3Xf
MBogAVVRY6lvUwi5w30Lv8ALM+HAzzEGuco/qRsLcRmYCUylNnSLJTr3SHmB3LQHQHoMRewsnclS
H69rZ2oht4y99H4uvK4sujcl+ZZNqlec4e4mjytdN/CxvF3JQ/rrCJEbqkDac0VAD3vtXQuQSLLW
4P1P0e01iVBa2FxnwaOboq0MFbdCBvmjcfh8GrGBE8hJdIF+YhuaRIWJUh2KBS4w7y/QJ1E1Rwtf
E12sPzH4Viv2Rb28ixOTDJBYdPI4tbZkvqTHwrjjN4hzGmAcGs4fSkNlErsc21LT2UYFj/wcpWO3
v2SFBt95p3NY9A4O2QKp18eXOLw30p97CuPsPf/8qNzWZkeYXhOZqyNFn2TkP2PMZGmGryPUSFGB
bMabhkgec9AaxI8y91XGcZ+f/gaNV8JJV25wWqlvBp824Ej2cHarXdZZp9h0UXvRxekoDCG9VL3w
jY886RUBltubqTL+1rsmdENH1ApGMjqpoaHH/g4k7/5CJelmpZRPdq3x4XYOIWME70ht7q0Mc4c9
3kMzzdF5rkIuUHGJ5ptLZ9RN2NsYjArNsLggMBIxBFiSBk1Jk5CR+IYVjYeQyw1L/5QtEC5F9OD9
KOsuF0zI3sSLCL3VuYwxLa3oH9Opfmp8oxUh7svruL5EsSftRO/EWTE12ThbzqKFr3cPTysvXDSk
Ag2A5JsPclF+Tg7UJizwBSwlLt1YByB48IcN7M4C95bUC4XUbL+eaX3utgw96XwFZRyfHlDBqHAd
jCPmEhu2ImPvNFdH5mCn1FwZdLbPgI4Fq5l5K9PqbHoeuDZahXdaDGibDVnA3uj+qsHcUq3ZPb7n
DmVA2UFCyDsiSk138VFrYUibF2aWYDTQYpGqrPMrVilWyX+Dwx4n5m9zLcbQqRdSHRtf1SWMNMmv
nbt+e8XABognqt7KtJa6uMnFRBd1G1VjR+LD80r73CTctnpKwitF+JZjEI8hgr3060bQtRTracww
tUpuOqcQe+A08np97kDys+H5TYlSmsgLHHjgP/uqSYw85WoFnyPpDE77HaNJxPNxWn3mEiCqtHWM
CO+vnGFWMArbAXNpTjIskDki2UG8vjl5OyUZ+t/5a2gRyMdDTYRj84eVlNuNgf66/0E7jgquj5tw
q23xtV3ozV25X7xm/pFuDWHWCYsTbcahx+O+lwl/ezN7ZuhJIDJ9gaEskllqROKpCebZmDf70rRA
jJDPI3u9iLkDN3expMEZ6bZ0+sLkEZhXNkeq9cKwLfCSaZyTYOoPH8Bp375MWhRL+jyVK5vaAIHg
BGJyKPJSAEiyeEAUHHOdLeKz6y/uKZYQpuxI5VUC1zBzwL+0ccnijDRGWUJxyf6bUVf42+wTXLyk
V2G6CbWDAFM2niJKtCxAJs9fC1y2KsaYOaY+uPUOFaldWo8kwIhZLb8PYpKyr6s+kLwl42fC16pE
TCOy/TWSPyuR8Fff1zBf4XtiHlfMWVbrtliJdzWc4kh9aUk3maNRqGmLixx4ApwsXV7oTl/gWGVv
Rgv4/1CABC5AkbyPdUma8EiLDSZ7n9fN0ai/si7eTHE6WqCLf3ScwcEqgs/vqj+MOic8VQ9eyKt5
AfvFZcvaPh7Ld4IkTA51D0ibeN0j+8sNbFWJrQAVo/Xu+83NLCAJIBi9mBXVBv+4xiPt6mOC5SBp
qiw+mbJmSFBThr0S+55eH9Z4gx4SsA705lp2zv+4eVkjDpb4br0f29PHOGC5HZyIF2WNBFa17Iyi
tVbqWF43T1F5L2KaAoryx/QporvoqSQzXOCaI0zC69vR0REo3lx1FGzNMkVgsnJwShH6qjtRGTWh
zfsEMjxqY2Ft2C60MASWe0P5PQXvOSXoykquOBi+ac5XPyMA6S30rWtH9yCXKNLwshNcWLTRm+oH
kEegdB8V3Hda02U3L3vk0m9mJuFuY9JXgl+wxLvG2zXIXmbLv4mOzjMcZffeEIoxG8IKcadbZg1q
lGpzH1RnkOjw4Jg1KywwHu/Qc9zk5c3zc6H6QW0xd20xfys/tcGXemQ5b/56ufV866sr9gfoP9F4
jsII2ojW19sAPCEvEuPYsNF4O0l9xOwyt7VDANtmunp3FETlglf7fHKV6Y+NS/gqIdELEXA0G3KP
U0QeRlsjsiwdMDrfaJ2nq8DcZXnsxGAzag+mc9zuBN3REU3xiYHS++DXnpFaiPLGc6ooVtnBgxSZ
M1TtsxmOKhUuAhpL87C0yLmfUxsoiSI5qs6qiTTgPzf1kE1GTmiM8P1gY3rAHnLtQ8DBaQRlIb04
nvG5/OpJhAev35yQf8cdYsf1mBsxMDEGPPTQ9eFMSndQ20pbCn2CD65iMwAvOCiTZjCkGZ2EuTNP
9YOpIkRznV53EHXlrxNHSWtbxfjDseWsEKP3IS+vhSvcVZNHJWi/ENOVojvjM+4DcMrOzg/iJ2te
JnxrfaYgdkUB7Qu1FVryeNO75oYUhHVTuimtcg1gSqrfN4SV48MDIhpXVn4aB1MUh6jRTXaTLGaE
sPo+GfRUbtKYzM2j04uLupsp8Hn2fl8W3/zuvZ/l08vt97NnnfhAIsTlqx5USYteIJdavZaDy+cy
0JUX/UFXyVHhPOXa/B5HHHT95357oFjckpOrREMRaLI2wB4oJZOX9jvzcH+PN37qo8C9K4SQUK4+
2PUhON6wQk65V1ARNL0WRXBf+VbpePlSxXKVWdnLmYw3bKQNZCKB0NfIhJ8JaXPuLI96NMLshQLp
7uh5lLjlZ8wfdYXTW1NeTsrHwZ+IxJG7STqUfuy7XqHvrAtc+a+k04U/gOTn5bToxK7o6LQq/Bfr
7h8Y9yJ/jjmdpoec3bnIllkh/KCpmnqjtCtz3Ct+Uo1CbPw8mI7YPSmb7jaUVlNDejv/D/NQ4FPl
jpKlmFo+HjdQEe3ybwdxD/bYIYQraSTaplGszXLpCFDWlZjlJWAawyknfVw8dMjBYBiG/H4Uf+oh
jUWY7NttDHltvw1JOQI5rzeikPKX4G2xFnS5DG4uk0Ea7eh/Q4HQrph4Fsn0PXBb0siHN0QHNasL
eDe+1HIIvsPjwjn1XPTB8MDCPA4++HhtYvr9entpp6oOUMbftKLgIt8vRPXzXpLCHaZMxd67VsiM
KETvndcUUwsUVwWjslBM9IqQZ+EahTlYSqWKfMS+RS0P/frtR2KiQcAityu0lyMq0mAw65VNU7xi
XzVG3zM4NK+r7cuNS7jMuQ10YoDKD5fI2DqAEvxZO2amA4bGtfY98PLyXe4jlzkgvxPmiV0f3lu2
fuFCmH4uCnn3pzVw8TlfN1pAgQeU/kQ19zb9BOSsHW4/FY8owkoE3RfAoARc3jmMi5Oe9rWoAayl
zkKdO8guItm6FmlD4MXTwjNh9I5hK7T+JMUl/mQ13DTOi2YWFvLERmTbg0wIeSM/4+LSBMBYjr2/
OG1JtTC/B1eDQZjdyZj1pzg0aIq7n3dJB5Vz8pzwCarVIgFYSMNbfueh75K8GhrKYacLKmBrKUH/
7DGEPLho73VQARTgY+4JvwS+ajA/ytCDRMVMxibGdccrzkRWHzXVABVw7YAHUR4AVgnu1efzWNX8
uHEeO5nDZUG4ZJbK8UPHeBc6fxW6udsCKP/WTscFIqNejc+Wc9rGqVoNk65+ZcHdgbs6UWNDTAVA
NYBI7JCKvqbWzAvEGoz+IXUVBTNdj7+KZUuPAd3lXIMnHsn7ihyqUBwUIjv4sS8TYpO1uxj1f6Zp
8xRvwK9o7kLN5EvnCgecXiPHsilldrZ3EXXaHLEBDYwuhzS0DHnRsTY7pPvxEMWdgMKynwwvghrn
/vPRARAmvmgOgyqNqp8MbR1G012+BELjwGN54P7C0XAzqLmog4bURatgchCn/ilb1HNWGZd/8d0x
undwWoLRPAlLPjSoSvi18lsAA1a+l+N56TvvqN4ELWLT8ihvt844Kdt21REWYWRvepWt3CFpi1ck
kBJoImCWvn0IQES8xIXA8z7HC58UAyahadA0x/BURSa6MDk/JF0LNlMbtLHVtf9HkyXQUD3FJluQ
Eo88aigWARimbSkgfwzwQSbEKrc9CEOPCL6B/HWg84y4/TgoxVW+vny665iboyoInTfW4XoaGNND
uSy1fADq9vuL8Y0lcT2Gpqhb/iFF+FLn35oLc1GEXU8sKvftANYloOqynOSR68Tp9VjE1g8gDayG
jgFxvTBp7VbR+Ul8lZj0n0aJhQLy07lGCd0kuG0JI2ddUz93c3oyZiimxzVxD++q0vHOxmqOb7Sn
KCguleC+r5TQbWO4atZjYdNYv6t/ElvZpwNfYoH6AkWjtYYWAdZiFbo5vGkrMnT4ttSM4IcP4w4a
caOV8E2HOFvsiG2cZHW5NL7E5JTdmnLw7a9KRApAkaBBokeFUCoSZdRn5oOuENrbE8LWKlDzofxO
nmA2JW8QqHfCFT6PExOcVfskLBgKv3pCuYY4lWPnGnGGVS5VGhzD8X8YWbfvvDFZxH88DSsfnnre
QEJz6IvDJjB6TD/aU/UqG2PYez/StnLRrRNhCop5haTzBsOq1hz8SI1jlrXNsm4vYz1wdPrnwJZs
UL3hOrxGYgJMum7MhVaZcazlfphhpTPpMHUi/8fskgMHQLZqi0fJ2mWYURO6/ic6yQO0D5ncwmjy
oSkz8JPrRQZr+bQ6Lp4d2lYZya2jG5veRfR+KxKsX2e2Tl6HHfdClm5/TmNcSbYkbQw07aHdPngK
3Kpf3LYmbcE8kx6J4Zn1Nru1u0H2kpz1dtMYx8aJacbjNLCs7GY87e2ZpNnEcsyuWK0PrbUtIKWI
9I08UlfXsUvNIv2b11KxvK6hL2znLRLhBeKYYiEA2/ky21Uza9Dyqyjidc2X2d488AZddsJULrgk
QpL2o9vV4JTTRx3Egb5DIMJsCmsnz/Q9fK4tGCPbpZQrS0hCgbkizPzJIoL4SoH+VgD1rfAW2AB7
WFw5Abfg7x1VgaSgOGvUHWyG4l4JWtR4cOiTfURn6CWwgJdE1SG70+G498cn7MgOyi8/EE+cTi7q
IOstTI4HwUGZ//qaT+WSk5hxTaLbKBbKayVvbn6tZoEhLMAVz2Ah7hlH2J9bm5Ps6Mf+vVyQRjl0
8apH3Ly+017xHERJGjUly/ysk68NBOt56bZe3coC1Cq7KkyIfdhOU2D6JaCaoxAy2X2QN6Iuz4ID
UJqVvL243DCSpjQt7c1In0jHNwffdlZgxIe9NIJ/zmV9PDf9aQGGillkCeMJ24fY17IdruZv9HJ2
6QseMnD10gUMccrU5rnBjk8D5RFGWGibo7VQaBA7QHOXKxvRPS/3qwDfyVe6ucCSBCZaWVFcm8VA
17mwjkIMwzyJV6zRz/ZsbsZPFVqdeXgjJqErQk+cPzmt1FpUBmEnAKmIoy6DTJ88YWOfhRC0CPaF
xHdbUjHIZqITUNy4m5Wu9+W3U9qwbgpetaNXmFItWCERxpVvhXyMdXtO97whJ0VVRCcuLLA4PWTP
vq1UQwpxi7CYRymzd5RmJeV8uvGavXRf0/V9rkiimZighFZ4zjBUp7qO59+dt7R71oA/KQFSBjy9
36kqw+1z+Disp1TBoROktIqfOS7xZ6rQhLkaUQ3+juWRGHzZhHizFZ4YpPVO/x4bIJrraOAfBkFu
Lm61cc9yd50o2Bdr0VpW7k9jEwu2gSD2rpKls0CKKjTBJlxKOXOXxv1erkRIBrh+QXhCG/8ssp+Z
wtNsNrJ7ymm7HO6m1ymkiDvJv1Yzhul0hcoV19XXat3JCR73bTaaSa1SUAhXUSGSl1Z3k7ynHytc
59u1F4QXAuJ/e/a+lWMw3CxWxTGKax9ZsOUd9SfzUbzRYK1hHLSeboXDd9/iCjshimDwjrX3pIm3
rTxLXrYzs+xkb31O2L8Cs4fjU5+swL+DP+hZxf5M87HyT+GYI8mrVSG5MmsuGuPUiXTmYy8/cLe0
ZDRKqgQxRyPNspwKEz732+BxI59deA7AAugv0iLZyZaPIgmga3G4anBDU5KGC5ztpqLhxUUabM/G
PRtEzArVeCQ4YZ2I5BCGfFLZ1m1jm9ZtoWT75zIrT4M1i/9f+JqO68220PbicpZK+3OoC/ochYx6
vjJHEF34rCdJZvsQ8iSdqAzx23rRf5z/abB4kqc+G8tR2HKINnghI6cuAaJ8YAyzRcKU8/dn4ruV
jdMwvq8lWZ9zwqvxpGUVSkmosWWvS/klgeHhCZM2oA/Y6Y6ubKzNKJrQ7W36FkOPSsE50rNcsW0y
xP15SgTvN/UWoDynoRB6VywkKQnSm3RxqQ8yIkHCw1xASZ0Na6a+ouIVyZ3/yuPif3cn9UPdtiN+
DNtKnlT4T7Yr1Fg+W3ylF8nz6EAU7OwHMhMDvdWuN5BY54xnLP6iYvYkoU+kJGBQ+vD31t7K8VIy
1KTQkoP347Ow/6pKWFHbV1GDvQU8Ig2b8CV8wGDE4kL4C/LJ2FJQsSem7/cuMoq4CnKJP5DAHCTK
jliQn4GObYY3gLBbHXUlquVrwVwXO7ajbaB55yEJhIAIN38Lk7kaG5dsGQ2HxV6GKorjjW0z0sPM
FvtR60Kio/InkCzSvP+elegieEABZ4KjAN6IRBJfSr3/WDB35Eh2WCntbs/D8o+lrPHBua2bX3Ed
ArOw1fDASEDuRXbGXHhUNTFMetEXknqLvZlgL1fBwg0F5xYuYBsMC3kpgxhhlvOUMEb28Zhg9jAe
pDUHQhYk7IG6Mvm8Q74Ed9yVNyQPcyuQaKdjb2Wtt4+5TWERTzcZdd8AsNvCQZmPQlpW8GSQB640
ZgorEusuTXoj+P+Tti3Oznplh+3imfdofbnv1N36EmNcuFimhIScVVkoRriqEoBWj4hOC/CFUccn
o8kqmiOAv4G033O4dA2Z95+oMX0VVoqx6LIXfY4Vz7iTnumKZEpAEso3Qn5rA+DmEe85JKB3xnoX
XVo6skYY9BbJS80MFYBYFhlMJ5GEBf3mqKgn4fUQoyeF54P23sQo29m+xIoavXjLuPUbYFlT2I7C
KjcPcyXOeQXD4VL1xvAPgI6/S49beUiIsLNMP9O4BtqVUjFmXop3fhJUCDp5eXw+0W6xjyAaDcd7
82u+y7CLFwXgnhZiLd2iquwnJJzD497dgb5f2clyM3p6RMaR2cT487anTClyN21rFWg8cWnSHnms
C4hcN6LAejaJ79V8XYSd7zJeTnp4FlZZzRDFeYXfmf9wNI5MylsSlTAZ2reo13t24ck34OeT9EfO
+/Q9oDpTY4fCtCLh+OCW7WY9Y94rQC6Utl8qvyIDI/b/ZkWWZefob226YrfGQrMJR7BVkme2fJhi
M31i4U29ylznRYPdX2O/GHqkYN/CQ6onZvNMBNTRDnjFCYWBKm4+zJHep9c+/nfOMvve2MPolfhC
GH2R9o4fBDc7s2kUp7HqLVVDzab1Ft0c016hYDVAMvb11gvOLGbhrjuG/aZLcojYWcUPTEaXLKxb
4spu7M9z7jbNwB77x+XNZwyp/P+l1KRWcrgjgghxn6RbDxOWzKrP6CRTSdn85mc9OT365x29MfT0
Vtgouk9ZyJpFmyEcQwZiNxAcv5hwb6NWTIIAgSY8G6+DpAOxYUIwavOGPZmDXbmdUrhX5YBueGr4
sGUsPksIvTlK5OGYZa6m7fewaSZ08xLv2Wzk2CcplMYHPst4/zU/gp9W/EU9/3TdJPh/qrGwbEA8
cdUurFbzWYAqO/BFTzp8YpRfbD9R5tSoNiYuG9muI3ewmOGs4ztehm4WkQrtYMDGA5jPNyKzDHjS
KyO/QjNk6yVyWYzE4kNGHIEVFHTUEVJF9/efWID7Oyb5QEqAtq2ndngEepGaK5RfJSyn7ue9hLF+
EDoOVZejo12pr0pr0wcoOrZBwjtehNIOny26/FIP44JlcO0U+WbrnIJ/Pj1Y5xggw9/9Or0bjkR7
jciLfg90E6flAfX75ounqmPCwDV7BRD3Ya8MEqZSBnAETqg458QL0yZetreFOHuBPR0Lfh6GBSZ7
uV9TOpn9JILOPVgsy+ZPpRXHiVTTS+Gkbc01477ev1BaZNV/yp4pS25RKOI2H3K/A6xhP95YIgE0
sZlmiMvPEvFQcc+P6rA3TfandSSNnkjb6Z2f0qm+xtEmxAkshe0Z+Z6b9kF1Z6UmRGhg4Oxa8bNn
TBYH7bu5xIoVTTTMqDooFx5e3rYjt4ekFbjMvyy7hW2l1VlPQ4OcBfXVGlVzYJcbi0VWTehi5Sgr
N8r/eh73PQ98kkj37EWHxk5RAvnNpDWSchJCWTb0mvXLkR2lhgEcUPRldU6rziJkx+iuT41PLD2x
MAI1gImNuKnGUHxwAAuW/qWhthCU4M/Wit2W3mjiyz1RUgENq0y12wLCFMy7NHuKhcWCgrNZQWtd
IztdPpDZ9JNEudRlfqEg5qvJoLeFo6I++HtVOOBJR9Bm4IfAExjq9UPFpbwun25aaB4ri09R1hYa
OBPRrAySDwjZ5o2KRTnwimc9wts7FZ12CugUFrqMDXo7rW4+S879Yj1ZN9Z3Yxz1UO0xaCvONh6Z
x3XIdAFOhHAirf9fvW2obMklBgX6F4YtBxkZz58AUhIEZ5jc1LkUw37EPbEXg8ukTT/FO7Dn2Rv5
vNtPRgxn9/M19o4o9wfZrqqaDCaBhmZZ7vnTAflfys+nsNhmFj9M4GBQmjL3E5nNiF9f2I/h7wpE
cv1grX4iERknS0AgcLuTU2Iy/nhz5oWCfR5YOiCcDuu7IN+dIhyB0nyWS/FmU0ZRLPiLFWHzCga5
AfEhTqvCqwdSWCfRiAmiGQdYKgUs754f8ij7MX8KbFfZFM7dvU0oxmp/gJi2ZtazBrwjrgOHc0i2
Gtw3U1tUUzf7ciN7G4Vantj4RylfCEiZRXAZO2HfBTtJWS7Cl8lMaulMP/nY4vqcvpOnvrLxKCFb
Ly0jUd4kqEUslfEQem+4RXW5VvtY3QSuGFbc/AnuWSdckYe49RkZ+OwU24f6cPvx7o18DQCpYnGo
vz17YlyyOHSYB2MK/LeB29LVAh5u0lAc+78GoE0esAZhEOrhUFraNIhqjpG7FNK0DwayLRS+mzMa
DYM9J5CY6BqGM74YhkRi/rN3gmbLV1zP2iuIUiOs4RckOIi+hNfWOjQZDWU/LmQJQ17hSHK/Xk3O
7vadlpeaSgvo1g4oUgdRdpwVHKBz7+K5h09gg84KYY83/q3T2h+xU+hKDYxLKdzkyKHg4E49vD05
WoDKnfRsjz900JRoxHtQhuz6pegY1acArZHNvrQft6BmFF5V3qdoLvlDo0Z2ptn9BU5qD/xw+vQk
QicGc6W5fAPLe/eHfkdxtlpvp4zAqWVgE3Or8A4dnfS6ISzSsydswY+8PiEoYX/zKaq+SBC6AIT6
eCWqp/4CMoVcdli3UnaHhFLvYD0mj01aC8UDlXgDeQMZemuINXwruuQsz8mwnbMlN9r7Y1Uo9B8u
IYzT+XJNl0LoqewGYctY+cHU/PboYetdUJySuNSFH8DaD1LhIYgAv8cRMvOPlcIguRru8sWqJECg
SmRMfIRHMW7kDs4jq+q1ht1vREoFWRJ9sawQ5luCry1QSCkEL+Hf0V0+ARCeYufpA356hg0L7Sii
3jpabTLsZe89UyMRM5t1SVtTpcsnlnNxm30wxggW7qjWCP/BROUM3MBYyR1AQVcrkYo/Xdf0EGS5
6q+0e42bIZj8DuWxRd54tI8572TB8RJXEJG4vwjQgSAMIIiASgvRz1AqBUzSuiXE6eg8pS4xIckh
HscrqgG3Kb8F1rdJiuzjg//ulpFV7yKnrwGnTlwJTPiZqX/BzVNZlN43MdLutLp0+sLqOzPgHoj3
WaHcBWelhkEuLwpPAtNbk2z9Z1BQnSLxhObWzCWDON5gmygJg2BxcvVjBPR3Zle8+EdI5mZp1gwu
J9l9WTtpUEeFjnaNk/GaG17Z/ifPz0XcwvrF7PH9RzF6aJQkuNPdAuH3Rw84abDGYi1OEY9kKs0a
URZqYVOS5IFK1zbp0LQFymyBkpxRQblu2/1TJyCPj8UrOPl/4x0x/AAhbKmscUWQrRDiUXEdeAeP
X4eexnI3kBSiTVhWbDKY5ZhxEJkgA3qHScKK2zLqNKiH0Kt/1r5IvWiI4wN0yNJ1emT805x09D4g
BILlgJzF6ll8D1+SYcEE8melLxpxWbBZi9YtDeLOVjotGrklCHZZVbzl3RzXnjk0AzddPR+VzUTy
ahEf2plRJPK9WvBbovYmN2+aTWdcdy98QSqOHO1+cR1OmoB+x9q8yPBmPZOVNSftgbDqJ8Xqc76Z
qLaXop/wt+9Mh3waM/8M6fmS4o46ABS9TDctnE01YEF0VphUGgYdCw1EOlKvxYHglER44v5IyOqP
vzOo4xBABoKAH3BRmGDx2h40BTvFuwpFZ81IuhKabmbC5EOghDAuynL+3ylhCf6kW4QyVgbN4w3F
cZfbpXA7fq79M0owLYT47gLvp8UPpGK6wMCQULBTfQQCD5fJnqUDao0wwnfddHJeKM8aZGor3VSR
DtK2d1SuxuNFEatUvQBbkciX6umayRkfheDY3UxBzi2EdkdP1LdGsxGNGgmPSLOJvtQrUH10yuzp
v+y7Eq30n8x7QDD6vDRjWdRmBDnyzeSbIxAswgS0TYN+LWUW1cOovkyqCQ6cFLQB/pVPGZQgXF4o
DHF4IZR114NWXHISKy4e2+4Tf2JwdSh3aCAtWTzeugJwxs4440M5MF6eVZa7gEcTS2g4B20O64SV
rk4GGd//d3bLEUMd8FZK619mRADDvG6UXGst2xd4Xk8gLbCImBX4AkpAJgxvx4eaKGvdwzL9dMSH
TyEWlmcP9cchenPpKAlbRII/hcdZdly9WWL91CPBmSpNsZuuwWf9VYChaG8fDGtT945hcfdWefgw
mJxHb0CrMF5b9EoJd1xpLQUUToaDJ6PhpGlHJjk1CBcBu5ELxcJmPChDgEG+ZgWlxQGAD8J6YmHC
Zj/2W9ibkFYsWm4C9bZB4WAXY9qCcYPvCI8qDiuGTZhkVwbI7YOz3OiVzZhxDZjFexVQw881k2IW
RVBglAgFkBSb3c3dYWJKkLaEUfHQdE9DkoaUhNuqmWw4zqnmde5ok/mJArFSbR56A3Qb2sijGSc/
iyEZu5eNcOtnZYpC/Mb44Jdfa23s4RZ0vXj7Rg55E9fqXZXcahsxY4DuCVw2XNVrj7xmb8xlx02D
ybAOnILwP2PcfblwDccafXD3Birod/cTigUJI0vEzs9rFzl+APDKqk8kg+od5WeYk/ZUnqO5bCFi
7RYDqHRgLi/CHB+pcDtP3EzQYFZKRMOSInmELoK8J/7gElebnc79X2r+R1UdTgdQWC6e/s34/iU2
XTBQImcunjb/VbEwsJmr1vvGixXzEwPMAkv1WAeVz6tckbS6O2xht6avs7DFWbDrbuKBRMJia6eI
/qsSK1guNZb5hafuxJ7ZCwQzd8q3cBLpaJ0mxfwhtbjudHz1PLcrBwz/azhIageMCYM0jFsgHurb
amuCq6cILtI0Q6m5yN8JRYrMxUAh3ZPWTs0JS1Zf+202uvd/PHUD7EG6rIAx/pIig4QP9RmTHJHs
7nrLCWWs9iKtDURmVdKcp7nhdFHc4fLzeiF6DGsSdfEL31phkWiyxRbG3TFo1SuK1NucyWP8RXWL
tqaCysDG8sPQYdJWlgxFbNRCSTsHG9hzV30uD752O72Alk1z18DSeeuIgZHIIpWQa9l8ZK181K4w
CqCrURY5S3AXaSP1/h2waceuioi1TBILEr2jwHnLY0n5Rp6SaFsuRU7BySPaxBbOuiWbs5GuJnuK
1onUss0a+6j1l+e/xAzHU7vntzooBpD/WSN/0ry20fpl5cf58t3Med03hGYPANl4B6NjY91yqML3
ZTm2/a0SRRpYHBPZMcZBlyz3Fi/ukAazUTw/vVrVTcaOcDiaFXITSrNa9toFvOa1Y+GAOMofpxDv
vB5pmjzZ/GBSvQDyerKA2Le3cnP0mqGP3HKvKl/U1zt+6oje1RAtAAqfXU7E0WvRtHJhQ3Evp8YK
H742s9UOu1x86wct/dpSxizEvDVKVTQqmR6ap8WLlxSRfhR0RgOBIYYKXlu+YwLPLtct6wO6AoYi
mddYkI+lIlhs7wmcX0aUJMnlEq/rbS+HNNb6GzAqEBK02FdMCVTRjpRFOLFpPVnWzQvApPpAO7rg
N1sRTgCmLhyTZsrXdW6eKsahyILh84jhU/3cNGAiow7QzoFU85EdgHujJ2L2c9hUH128CTIcUJxe
DMQ2yEA9qP3h49czucITFV8cglpFR5pzCXB+DvoOZLVhvMxktPYoKJSJD5Az6wilvSQkkaQZR1iO
zCybOphZ/HZBnEvSDvQMVw9nd0xe7DVEem334oqv04LCUE5nBHD3mcMh819xeVmsM2nEdZrGSCgI
Xq7fnELb6RFwIsqPE1Mlzb+9HnkhV3+cESzLKrl/Dn+FpJlDNgEwBtKXodInxml4pznr+VKN4giO
1P6BRH+0llwSVz/7WkT2ZlB09rL8cYo4iyV0L4KPFOzbiGKGMa2ioPqF4kFBQgfZHf5m+bfaqXB3
GTEsuaIy00Rw6b1siwXBg6Wf1rhw8Rnkixmge0URY5pglAtdItyL9Bil3altN8USJIb6p7u4RedF
EAyQ3fK8L0a1Znves9BsstwQUeyEpG5Gsn4CyLq3hpVn/U0+jM0DRWPGQf8zSw2s2wuNF9ZNrDll
BxPKipOEdzpPW5Rr6eW5R2pRbpQt9mtRXVsiHc5q1RUXibNG1UAJtORZGQfBJaaCKk+m+qjrfmp5
T86d4gnzBaUw46AeLplJ+ZAa0ly53TZ/cUCRCie4MW93Xltj2pHx7z8Zs7in9OjZpNMJTZN4pNVN
16YwRhTjCokf2/upa7aXotQP9HAKHKSzvsHrgYtHJ31wINTqvSHETka3ECkaexWCukgXKnUNEOwo
7c1otdNLOtW930XzxSPxHWO9A1mFiroYHOPZsrxnmyaBI9yc5We1tfrzZsdgiveIHhjNs3EvXCC0
6MJLYSYkYG6ZkDukBMduZ08gzhwX30m0fZdzjATCgYUCGhusaCXWNnqucYQfO0NEJqlTwTPC4hNI
qnCcd0rXMiaVuwOT3V1Y4a3vChox7c/j9Fi/TDkVyEGI1nGun8CVmX4YIBvidgM/KFFRfomPvyI7
Ki5vSUTH2PoJWPi+y3jPD9V3UnlCu5iSbQKhw37hOMF2k1TSedv52kHbDJfni9+H/1pGENm3+SZN
P+SenTijzm3fq+iaWqWi/ZGYs7Dja/IIhRS60hS0RlIihaFu3OuGW7I+CFYBI5OLAkeBRI/7lv8h
vr7rPw7EIXOIFlXeHAFZTh2w4MzXBRu4Wz8l0iAccv5DVNgPN6mKjGF2btmpklXlE4dUWU25dZNJ
oz7JgmCqKa/REbgdNkkLgLQ6h74fe8unhHv6aytChJv9VlaPrJYJhINbsFWsj/Pvs0ck96YfRfAE
wvbjFAahcaUQpeXDod1zJW9/DtltdEXxgw/K1U8q/fNSFOIYv+KfF7pWhW7R0pAAwHc37PwKfVMP
6CqVaj1apPEAzJ1cGPMCTKkOAtzsOTCefeHPZTj+mTuibeZ5yxmgQpjX6wmT+Ex23Ci4B/2eRHZb
q9Us4jrf79JxVHKGVSVS9JKUoYoOGxlJhFiF+7A5C38+rbvSZ1VPorlUIaCsVC7zBo5Y5vF/F3xR
gVpWezAYJPtbiSRUDS0pjnvvwGPDLq8ZXr6PVPQ/ijBfjNR5ROAUqcXt2IGd26d3ZA2XU9nWOmP5
BSDnhP2i5vhhXD5BwoXB4lDnmXaL4WQ0PuSSzOuRwsJzFngvqgcgHE3Ywc41ytOTaHr+NFiigk1+
/4DvTLHs4jIyw3gNIECP+bXcJvhr3lMf4lznoIMuJRvIBDas477ZKBtfktA5N/u1VlGuY6Z5wAbQ
s2UzC37JHRxx2tVbJWiwITxNNGo/y9MV4iYyDaRDAttTADMpBXubXmO8RS6V6rA5C4rUe/cFgJ9L
dRoPZBJlDkXWLpEe3wFPxHDc6RQKfWHekDokInpLUvHVFttR5bu87K1o64JNSQD5A3Opb+SqRXbA
S/BDtlbos6GSOa7dwf0S4+FpSagvjEg9d22O5s5EATeKQ+8m36YZlPuD72vp2/vFCqcINjLnxnTz
S++M9JoslU7nYfTTG0Hl9uW6ReiUm9bpguvHcT/y2OUQb4dZFbvXL38vmdtH5CEjJE5Nwd+K770D
7WK7vIiOROC7uwo7lkrx2oSYtaQqEZqJYPw5xHQAdTTKCtCwRBzIc1Rz/9Zx+Yg6MW8MF1tuMQjz
grBZarXpqYcYcSUsG8/RnHU9AyVbX00m3WdY29hBRr04Ll4xblbJQV9QCUmMVMAtGGPJnB01jWWx
6ecSSR+ef3JVz6MOdTYc8R4g9laF5XPWf/Y8lgk24o4+ZTGihCsX8G9p2ga3BPKGQCqR1XW/HL6x
55VQM6c4dSbTJ2UsNMPsklC9235CGgc0UYYavjakntm4J/MtYHHUPw1s/cQMDucjdskuAimg1bV4
fy+ZmufCM5oMpm4zQTgjxSOBG1agCPva9K0SFUFHlgbRnWkL/v0Y1CCAmJsxG6lIc4+6nBsroCSq
cttm/RSf5LkBC6ZF8FhOBSJyeFJo3fM0NOrmWkhlSK1zBpqcDf4fKshvKC9o4Hu9UoTauyEJyJja
GHuLvMBP/fv88Sl3NIncu1t6+XuYOwikrcGMf1mxPDG+4V7wBnDnkiudwmIUluF6AnHjlaJiJQMn
YAXqv8P5F0EOnsk0hacqeffzO8BkHdlywdJnbQ9euFasY0GZkAbfzP30siPBLXBrT+1ncIxobNpt
/ubylfjVtaryxLqONKuBvyBMfttJedHtGrZq8MWtn5UmZYsxtPKd6inu3eMqvbkiy7POinaTjAH9
D7ffnXbiTSeIFbVGnB1yS6ig4CvMrlPoVcwokXPtoZCfSvwvSYC4mgsxmxqpCq96N80xI7hRoTmv
2mBXZpchsZJ7krst4a8LQ0WwKwIn5PDaVrHQIaxPxs94kUmk/5UzIBTxcVmE9H4OhsiWJi4F3FBk
7hIazwqatIVdqBymXDicfv2Da26Ix3+Oq2W8R1oNEMM2sIDpuu2LYE9yyimhuA+mYwL2z9/W2fZC
yWjsS5mBF/0vHx4/CmwfgjigGVTyN+JuN6GXoODp2G74+GGN7yOGLxDo9BAqC0Rxi9YDVNpHkzZ0
ZhlFq/bagszikVBWe0JQApfR7Oo+ZoXDfxR/DC7/RrF/fLhI1jeKngFxcCoxL1S7iYz5j6cIdz3a
DiP9ONjon1iWk9qp4S6CIKGDiAPa5YghIAs9Mp1Bgs1ocEmCfWT22zacbPrtcV12HLgBGEVhNXt+
wzHfvy6DyDW9POOXytxwdM8Q9MGfUPPho5kdcZS3/LM/jd/NwqnkaIJqm/1FQJ8XkEzzuL4xWpzr
MWB8dGHjfnMaBgnQ7vQDcvHNhPZLz5Hy3n/bbC7tndARi3cYFDVdrMoFVRhR+s5RrhgmrZ7bqeR0
KwlhiHNg7nR2q4zyMgFr9P2afqZMP7ynbwNE0++7QUiz6BAVf8eoc9pOqQR7WBtEJjssKa2nBCb4
VqTbU600msyx2FlrObjZyvwqaOLoGGAzkDl18O4LNo/zIMaiQZm3vv7Rj+3xUFxb6nwuHGqQ5s5T
alN5uD+3DY5l+yd3qVKA7MaXDiDEz0xXm0EbC5S8nrkCJSnOgaqdVKXWQ1Hq1aCmX5CYfEMLB3MM
JW2tLI9p6XimdiR3eTP1BKffrSgkE75HV4368dmHoDvGf2Fq4S0ojCJfzcxAAKjgHxD3x5S61fLA
TDVigsOLAsxv9zXF/+5rqHUeHnU0fqgY+ZE+Pq16DZUgHNVyc0FIUjGt3e/rB07sUQbYjD/H4UM5
eyUqJGLnxAzVGxQQc9aYJtY1yxy1IALk1FvehW68S6FR2Rd1pAj5OVi6mHfB13KIQ3Q2BkRh6DOr
TKKLoELVCc2sCpddiURIzr2hZZMexD0QT5xec6fYHVEKyYxJ3Nr7nxm3E5uDFqoXdWvG5yTO+bSr
LzaCdWssRij8ZayFcuTVGBG5rkqyDqXAlROVP/KTTZYgbb+MJMK55kqLB6BtqQu0wXb8ld/BYqOt
P7/x1+c+TURxgAWuKdb48DzynU85ylHCgNc5fKh8ybqzlt63E+mr0bUwEyeZsDlPEts4kO9+yxmR
jBAQ1yvcExqtT2GEP3zLxMLzIGTZyV+mpMDRLQlg4d1S6fltV4FQWTFuiaGq3BdvHp9JU0c/PULC
PvTTJxsQjvi0mbAJU14tcEMJDEXIAxH8PuHAmHyvUH78EV48nfKhtUmR0cwznjRJfrWYXUhwAoF9
DNEcV2lAvi8XGXBzHKfrGhSpkhgr2c5+Roa01nVPZDyq21ItY9hoovAWxyumn42fLo7FphRML6T2
WezhJKsl5IhrQyHggYJEOECKfltaBSRKn4+W4QiFRXG432D4E/ceROLbIWNf5fwvgrXvSgup6yl7
XYuV/dVeNKLGrw224Q97A37zPw8eEDNkHc65zPmsTFFm4EPjkcLN89yXvs2CuUjMJWYoS1jDXCjU
EZDogP6YTKgW7I1n8hqXa/azhRG2P/Ubob8nMuLShbyJCsmgtQxgrsuLp4GCJTLjrjilvB6tGZE6
hZqV/iCxD+l/e0nLCcYTGe1QhSbinG/86DiGjmTge4Ci9SUAloCRv3dGKw3WkSqcyLG+Z14r4XFI
QUqOoExNvEvGnjdhDDqgC6fcQ9TTSUyZ1W8VuvWYJLoYhWWYOonuTDB4w3xUP8ipvqYZGx4w83tB
SZ/wqYx4CjNwGSPXjeSiE6TnUQ2CLwhlP0QtmsgpeAoUTpMUMPYDPOKxwiSr4emInwI8WvmePGvz
z4aaVgb7bTk6IPppgS9D0jcMaqWYIwRI62qyf7AKOWDpBmJF2JKH72aI++TJ+JXWFViJjHMpIQGl
f0xmhT3bQW2S2kj8cw53tm66kqPcFl1c2uGuTuIwumby252LwcuxP7DLv3/taLA1t7Ef4zqj6Pyn
g+6g8fHuBAYIt00YTYvfQd27pmgbWcX33ABo7e84G1qmQ0qiuqI89GQti8Ck+6kjnP9DcNZjJwCM
OjPCxQ6HMRSQ/oAWcSaUkDaL1oC4tXpqgYHvj7p+XeyrL4YUBwBLGnS4atk+kY7+AP8pNxlupYbO
vaR9SqFqJeEHWyeyTazt7y+sPOkioJiQr4siZBDcXm0LgAJMZONyZ3APtOgPc+lXysesL1NxX6Il
JCcb/Z65isJ3RoGuj2NG4UAhGb+660/5g8/Y5vkqE3LigONagxLeC46BO5JoMNSe05+EtqLqPq6S
x/EZXrNLQAdlpxKhrEqYpfUKTi68vTYwaphjM8oPbwZoOTw7jtrsnjTwfShTi0HG6v8XIvFK3/B3
HdMpf1DMKVk8Gv6TDPrt3uB3lZ+LPXn9r2ORlTnq8acijFDRMaIFNv+iBRIx/8eKHk79l2eHrBAF
Qnea8Yky8WQlgFwXx+7goD5Zz3jTITdjtHkhQ95Tvv7Uqesu6krgaYO/XLFnaLSMIxfCGGkGBHG5
0Et1OoK6aBG8mzAGLxeoxf6NOd4ae5Sou/R+bzeYQaWJg8gYwWtESMJYZa/QM+YWoCy799TDaheV
mYDUmHaT1q78P6mkSxdmyfAvJdbFvuYoRREPpM9PbpSw3qSnhf+19EHWTbSAD9ogL3uCV4UgCLYp
NhU/7MPt6XF5cQ24DBQrEqeCPcLbTZoNeKtKTARN0WKg8Ww8yLkWSs2xFMPEKEDKWJPYAPfpINd/
W+msoztelodvxns7m+xka0hwVIE9aAgTIknyLqV5KBJ1Nmjka/nq808X3M1hy5dsAuxAWUPkiSOu
BfcL6KEcezhuB4QRHoZAWO2DYLriieh12JqGbR+MArr3Yy1YBldy8KqA73hAptp/WK1aBsJPuuxF
OZK1yx7F7y0kuemR5oAoxXYul3cIi3tL7IktT6C1uuNGuiVrTjSsvNILQfMrMdF1VeHxDWtQKFca
zBaD8u9xhYIi3VPTo/tJIH2GRNWOKBnfAbKQH3NAhSbUat7bj00R9TDnSbEM+uCxyOtJXiT6dZs+
M9UD7kx8cI/1qaYzDinK10moUtvxEQsN1tGyysFFHqTs0/b27R5nqwuHi53RMkhx0bmW581egdKN
3zS6PVyVulmtGUEi5tz1zRUvsK9agWd8qq3XzpxEkuUVEIao/rao+xHchM4egZ3tyrqZ0YcNnPtG
+KCJP0jadzH2F7wVIM5JB41rFlEoo+CyjeiitKirIqyMy1o/34Wf9SKZ8uuFhdpslPbd2rqUIolC
Jfss+Eh5FjdOkrhBPqadjHa4Tmidn6uyJ2MG09JURoYwIgcmPvQbQAztxkUpvjEgg+jAVldAMFQ0
CwCuMSkx4ykIz+izTa+m3YsYqkFF1RpDIe+Gx6tj/3jXo3qtDFWweNfZTganpMfoDIa2Cu7SI+hP
98Pk8tpzYxPGh8GUQFqW4HD/yC26gFYd0mybXOktnZpa2EyRbd2LGfpyxKVGOy1pqtbxyOfCz/NK
hZii2HR8q/niiu/puGjBA5z3GQ7KjwTKfQVbspm7lXF6KAfE1sUZpGV6aGWkHfd6EaXB5bVyg2c3
qrdG11DBjhZKLIbiVTNNRZu5Khf3yLOawQmAQRJOH4LPfQoYDagomx8BX3CbxjbnM2GUwncQOy6k
nyQHPNPjt5lCjIDAp/AxbOqwTL6IZ5B0xfX+8Mx4FhhKsZlH+I6L14mG90XoHyW1p0n78GkABGVv
Q8IsKMLFjJFCtmjUC4pSuRLC8AQSs7Mnk/KsbRfUZ3FuynLT7vap1RCoMTajLxX2NdVzsJNdMKfj
nNfv9v9zMrzT2ZgNZhc8KFReufBUEcPKnydylsRx46rd3zQKqspGDtTMai5fHTc/UywJpvHhuYB4
lTSfEV7EHY1aufPJy3BXUHpv8AW0i49mIP7JwGIAxgcQ2T14lHErhzzRQ+t6I0g6EnH0FIXo2e2E
ZhstrH2KBu0gt3tSMYmN5j0tdrRxGxU0WMyy4rbPe4ASwF13RGeJRoaQ+01M8hS2ywFWrko330eH
nBNYB3xplcPcybYwQ7TPRx/mW2Sn1DRlnrz7YQKImyqi+xCbHJypVj2zHjL1lWZ8MUsyu48QzLVY
j+YF26JgmpnkejwDN5TllMCzgxQIsNWfQH+7zeysmhL9onjO8vnNp/lxDxadKekpxoBlo3idGjIc
2Bj7cnKZURutcBH4MGrz6utqIfWKwH03bu0LGQ0JayR9b7BAHidijHRdKCnttgUNR9o1amDUurOL
5b9YJN0Sb3rcamo1BrJLVUbsG2lv+Ro2woAmP8gi4DMhgl5zXZCkONKxJ30fmgN2KLMuzmVguBm6
hdwUhDus4J4V22t6uzLBDlMgCLQ4+nOWFCyxk4jx02ilBbrXb0nXoI+m8xnmBKHXKPlDZBZh0SEO
XbiGL3g16bSOwat9dTnEXG+HNfER/0kpq31RC7x1g/IHGddRNhVpnQ3fOSeJGZo/BBXYbTsnnH3k
dqKJQI2Du3AgulvC5lgfIA5AI3pa/E9qvmctLwkqzWOUS2ZxF4NntLBrNqFlilQK68jCXz06xLqv
b/0ilaFRqOVWncmcnsFgXGNArBoe7edm+q+yi3aKtCZ0iRaUTvrkL3f7bkEyHTzZY5lmILFuU27V
nqgLFod584tUszsd0ZN4TeVDYS565Lt0tZEge0jCS1mz1kXrmTT9YxgVK2IV6YvdB/egv6pgXis8
gbBif1sxNbDDyvq9Pdr/j6zJg+LJX7ANKtJitn0900pe0l++hdnrlkBjvMU37pzF8GoXJUoho3Y+
a8c+mkcQKA5x03zt+qwpGnkGUyL3cIea6yP3+aSFxQil5BRUhGrWRpTmQ5phkC3137HUuB0+PGE7
nX6g9WKQ2WhQiVDocq4mYU4ZbtWEV63HusQv9VIS+OPR21T5xul+fiHO/1T6/zKUBqom8EyLwQUX
csHyBPxFbd4Jb1xVZ0mBjOsOQ7mmgKvW4Ny2jV3ggzp/dEaBMj4WcedM0rsc7bycnZyPDhUaQ8Z3
YP0irXsY/CekAsRBl6dEZ8ttmpf5UmnKh2/6zvLjwzCDtdC6Es8Morxb2cyTH9mRHbnxcTEld/HW
2u8Sag4o1sBmeyrCWRbujo2EBQ3fmCOxe4b5GkN5gJdR52w6ETbspkHDLBX3dziS/9UirQmyTrlx
UXPU3LxkwMU1UEaqRbFPirKLKN5dGEzFoqe1KA2HgOHBpaJIlWYn+4TWvPgfCJjDyJCI8MxhORvf
w0GJr+4KPLgjYdccC5RrvW/3NhyQamlgAgqfjmbn93+rHkQ++ciF5vTcLcZwUsR6mQyD2MFWKkWl
YpvVRKT+mL88QDqx2NJ9qNg8Ded6SIYks9tctfV4CpAXSnyhqfUEzoj63bYaS7xhZ7L4PLXUS5Fu
y9yhnl6znsiWwoH2jZqenvPkWzF9VCEbt8W11SlXhOWYqNZcl3A9TbRz937zE4xtpQswsACmpdbT
2OrVRlyWP5bK/px9BaLN5MI67oydb+tP1gMgGVdAWP6hjkPHGishqocIdorJzkp47ZeRFZdCvmv/
TKW5SM+39XzDKvf6fXSXRmaCI9pelTmpG/fD/a3KI1rX5cGwNEYQeSSnl212T2wFxnKSKvuvbtYU
RMMwH2oX2iQ28yviIO8kTx0w7bk4A4yHxaZQpt9EoUSJ5j0TVbu4Kp/QB6xxlfXCnMGm1xU+1fJX
dq00sAPyQn4oL1jQoWDCB/1R5K9XWxHDqfnpofPlgSn6toHQs7vzQ0WiDalT5KFCnLnuUTGB7Dnj
4RmEprtCqFH9UoSORm7CdjZFggj+Ovk+TJKIOLdef0mhUxbGQgRFEwo2oq/E4u2z6880Jefw1ynG
pfFxh9fwviPhOiL07Tm0UFoUfu51oUdPsglCX3uQTuZ0BWUu10nM+Srxf4vyPeBnjK9F4Lc+kovR
lv5KCgivYUoaKZBVoo4WD7bNmAE69KD7j/D66djXGdtIhJt5U2+cTCvLoK6N9gCbbgrMy6pD4Zyo
duV7UBgam/AErP0CKsOmNgiMM6MD6HuuyV1UOBSNGxPBy++RpXWxGkCSAOpWcx39Tv0ISug8u8pd
QHs4yatAL5nYZrOP4GpIR1FKaFMDKn8g7BQPmLJeh8jwpSHce/q5J1GczD8G4/GnFXkeEv6mVQeE
bvVdoIE9XUALOoKGdU1V7sCoBXIz2f4b49lhr0gNNdTesuZ92PLrWC2do7iWsxyWC0FWRUUSq3UX
OxjpvDrsyU8Hhz1rsP1Y804BAimIu03aeWelYNqesRQvTmW733OpA/kjNC+HkgeMR5kH7bnslMqp
FgLTVNBIzxpb32afMfDWY+9qiV1Mohtf8G1P/sgeXR52e2wSX7tdPbV1tDIDA1c1eFn/cbsW8OCD
OzONpNIImEU6GXmKyTAIE5wmMBGXOPss/Kb8BmTIpKte0Cl310X8Kyq8SclD8eiIjdIlnuOnb/i2
vJgNBNteUw8nNr3hgVfqsOIpA3qeZPgzd0rb/lkAHCq8Xn4qKK2KMZsHaYqyozbZojQSQf8HIKiI
eCOXaFnoOYhgKy/PH857I6uHeT+/IMzUS7OLADwh5daTVsq1WlOKTaDA+s29f2+dWpLgu9xVT5jq
+B5UsBFf+OJvYYedWX3lpX8nFJroW5VM6a8uxOqQ9YSeR84nGShPhz+AMsY+p/AGfcgzHclLJi11
V6An7lF9IIRj4O/EBvdQcLXEmJi4BtPLzhv13OdiwiJprd9OkFpOQO0Fq6qeFa0IdaMUa7oZitKy
+YzgvaPHmzZFrKrtfVOj2o6VMSd4YIDEhtFEdV3Xm5iaL2vucIf6GEC7bSzrj0pse9gmkJgjZ7bO
1ziqxhfTm9v1YNPzJaeYsZq0yp8nkPKDaJP/Gt4RFIiNijzNn42jinXwM4qTVlfRK8/HfuFpHl4P
+UpUJhFTXrTogBP7V2+dfS6fn/mOw/8mRj/05bdo/vccQ9i4xLeUU+332I26Bu8JOfP679i3Vss2
kEYiwC24DjGUK9lU18Z7iivs21jcb1dY8U42DckVj/lQM249DJY81COZVzw7LsZOhMFhNxxYJKTS
LuCkGKce9WtS0npiywOi6U+bGUBBYwA8DGBJWB8NfDPYv3p/50b8E7v3B/Gzk8RtE+3/8DchRHX+
vh4wMqpVISLZw0VcJ97O6UdixzoEedGytjHDHDiDXwtqD2NkBYGcxQoz6ZyZeL4dK+9305QPSPRq
GSEmfXfF+/eJB9mTqRr95JNQAgasvbidFT79QXowShdE6CTFixT8oQhUWqHqq+G9PwSl73pNbXWT
ZBu+ycV04aoCHUTObCWuYCKWRrOl2EDPxI+xHW24KDWPb5vJh54Fyk7mVjigWpIHQQRD7nT+Q5jo
SWYTJN32LS+9Z0sIEZiJ4zUU2g75x3IoyEzNZfX9Mi1A4y1BPSSoEYGBT8CJx8MypuYfiQyT8dFp
tjSfTYwxG5u8auVM9b5R9ESzRSyVSQRUGE1JXWMfrG4DdFWJgWhF7LvIgq3L2CoQUSj6Ncy2yHQR
PwtU57i1n3jb8BwTQ3j7s0nR79TewBTzFw/vrZ4l45t3vbbPMHoAJ8mIJU1+zDgfakYJhggfK8kg
83c50aq4Umml2I1F9o9wssDcawq4KD8WyOgfNTE4GEsNLvR+sR1NNI7y42s539PmGFsWczaIf6lo
m6h+yVwRucKaH9BHtEOnYmrqxF1xoFgOi6OppE6iv0oqRM8dKnLvWDxdhtkTcPaybrK/DxMAwgND
9EM9e29t/eswB6YlMBjj8nfcNHBldj98jUOyhioR6U51h+Q6dVR7zIjz73dzrpnjN07QZsj1vfdS
xk3hGYPJtKN+M0I1s0kkVW4GbV6qaeFGvZW0zhZAqsQhMkfhu91VfyX1BJpiUzHlrdQoYY2VwaM8
TP711qRt2pfpUhJvr9z0Tx5SbphAadKdmlHrP1aXg9/ljbFqAX6w/j1AcpD+Bxjre4pd0Kv8c8su
Esvq894gri71SOdcJ0lcl78POCPNSLMX0LYDsIw7nNaIQ8eHwurILhYKXBUBsx1PcsO9rwX3pELC
FYoMnmkwH0kSO+mgGMn5qIvQSkXyxXpaD0mF2Sd3KncSIHPU8XZW4Xz2C9MiIqdpPBNVk5tIIA1Z
UVB0VBBsGXSpScFXxCX6WJn4lkErMIcjmdUqyQI4yB5/Jz3234wc+NlID/S1fphDQzmHjND/MHoy
Ra/lTdK6PWdlyNe10a5juhkyvX5WNpSfPse4xl8jJ/rAjj1vicU967iDDWunJ+tvHikCzhZqWN6e
FL4XVht40vHQHpNl1CT3OeyrEpL8FJ1YmJiRVghssLYqDdfUxgYcg5e/8NRHEwDn+yb9ym39dBNu
lcZdKrVeWfJEAQ4Ur8XCDVsX8J6dM5TNRBP543jGQ8Y7RC2QGJCfTevpyAlM8qGFteE6MVuncxFI
aL2uJVntmGbidq56soqNIjoec9CjSqO/erVFPVO+L41lOXQdwT7Ssi9xX0R+btdPnUtYGb7mpsrg
bGALF48jbWnzCvIH83Hrdr9aMPcMAlNWY80RnMeVAuJgMWFxTiL84ciIJPs9i+vwJddJcF8ffH5U
yS35lCaSbuQZve52u0DJ4uSlYSCcMBS6ndccgo9U5HndKGY6m3kJI+/7/Atr3tL8OxchOstFjESK
KMgvh76erZsorakOavi5g8KN1NzMcGsgUAWRgP00UET2XnGqTXovQlHOlUpOgTQM7kIAviU8y8sA
jYpEy14fktnzAPI0PQYn3eVCRRH+HSN0wXARTyi/T1AsWTWo4mTB8YX27704gA4BRiGyobpsz2ZE
wiLFQUZwTmcoh92blC/0UYpTXgYDscX4EjWUb7NxTE0IWrS8/6FOyW3gUaw7OCbj3FKexFYYSs1V
rnwzu6wT+gO0Ws9GwIFREnrcS/hu+JRHJNBrn6ZN18eTsRnu4dMnZAKcaF5YFxI1NRzxSrCf+dYB
uQa1QUgD3f3Mk1tBoVLFEurhdYwu8lwGmb2Emrx7Exma5JqUaHk07nXu+ZqsqpM5+DL8Q6x6s0+R
RC6biZufjrobzL6mcDFtOf4mf8B/n3HDYgCV/IxMTj1RoTsW1zhiGxsunakw3g4oU2DfXjSzaae8
2kUpuHmib5Jyvk7d2gg47lzi0rsEipBscHleCWLNxSO4DsvpljN7Zzxdk+ltVM0c63W756fuH8Av
L0xJZ6WPkdPIIq25CgpUeVySPJUJ51lpk/kYBxYWVsL1hLpPRCkokv98BLN8Q8kF2tkK/BfkQiOD
k70Y1n+58VolHTZ05mVQvwF/n8x9lwPuwBW9BNq2sW1WKeh8RAfYdUkgcq7sZtI74Eexi5p4kB1S
FJL0tHkRqlIHbnHlT2D3z3Q6lpab9w9wEt8IuHDcM+4tt6DOUevd7rFez7Fj+NHtjyz5YaPKebO0
XnbP447E8eEYpq9wKWxTMd9iuaeWuncq+alrSPlDbBnZnRDlwAUTye3hRcxpYQRLbqEhyFnfye7O
po4v98VgGbEThI/y0HiS5jPed1UTru0Gc/vIKMx2icMKnBF8fp7uKXycrGlwFfi/k0jxaRWozMKb
49vXDpSmNZxWxVVenKIilDI6ZF5+enyneu9gWVPgR4PUuUTVp2GTsy442GzPqHnCwq8eCMiGMiCd
Gv4y0o8NvZnWGJoeTXUp7mMTiyohZk4cvoFssRi6QbwwY2IVCOa3ZXaMtYg29TQVvAMphVixTiRx
vetYS3+915bf5hy7tEi3esrVgOwPCdjfiaBD80R0qewAIhrXef8pctu6SIGOcDKYmcW7Rt1/h2YW
k2+uJbCwFI7JMfgG/pTSgW1NR2DeGSjFq2NvR1vEkfdMgNGk2fnc98Xkt2n2fQuAMjqesM11Y860
oTUOxl7TZw3l73SnN5m6Sfb+2/O5Fc7rKgNu1fV8AlD54NLTs5tWbC4z7wW6s5HJcLKqMpwZ/Pil
QhGfZOyLspPw0EswI650oKsTaM36fSSDCYSlg9mW6XzLenR6nyouw/W+D2eSfo00H9MBB9EhzUiD
KxG6vyVSQnIhNCnHhZGJh23dysa5sItQ0cv+PJCpbphCJmGiPwDHQML9f42XpIAecb0wL9ovRPjL
oTI+wddi8ODj8bunI4RMI21mc/I2I9iqfqF+qvN1rLRzO+TrTgSlUPevmGUCKF3TCqiNeGtjfUCS
9OLk/Tm+hK9ivI7o8hqJWLJHSs9tjoWpsRWjkjaR1Aq2hmGRwo+WtBUfSBtn1kZ7V8t4uDWzxRv2
KNrXLAjMIKWYbW9Qzw6HpueacEfmhXUqYMALb6hbBMrMFRQwglrNkpHG1/N/XuihmTFnq3VYw2qu
5qlh3vFNBqqgcq4lLwK4KhycA7xsLXPRLGYz2O4QW480XbDm8Ih4H/vV2ZHzZY7Ts6l6TfbISbB+
maxC06cDuL3GYWPMAU68y8YK9EiuUQ3/nvD95+AOXXDJ9PCW62yVtZI9uO+miTCrk66qvqRcGdps
ZDsarxiku6O6QYG39SiNn/slBZQx5Vx8wlJ2aJXI3bk1Pn/+fORlgO7vdhFJtFq36dPlipeuttAE
5j07e0yNpju4BehGFXJ8bvFKylaI3V5m4JDc+447SwOs0fB3IwfkCnRUnK2k37FxxJzQXY6gFYV/
TQc58EF8d6J6LUiC/79zQpmjrU/WD4LRVHLgZXvXECZXafgeXvkf8sjHoe6rkDxq/rS+2cZ0THG3
W9Xf9h6IeiRQEnky/2aN8M69gQtA2pZZvSNXv31o4/lXktaGx1Tx8TPYDAFY6ce2MZD4X2stMTbO
iaTz9r8loUizwzQeGee1Ap9g5LfVxLB3FF91W2Y0rAwTKPWjCC8YpXaUCcKxTbFTkQKHQO3SZmpw
L+AO5cNA+5K2p+NHaNH8WvSBOG1C3JNH/AvndmodGIYdjyk/UEJGVmK2Zul2nZidMdk5nYZHmzLb
SMiBuLlenBB1xrrlJWBZiPApocrQ1mZ2as+XpNAT40vkXqFr3Kn4WJjTtTQZkzUa3/hRG+5gxeqp
2BodpswOwby3u6UtZa46VlScN6na894BnhUJWAHO1gvoxXb40f/qKvHmGvgAw0XO2B3nwl7RS6V1
JL1dZ/CQT8fB0VRReGHyynDGF1RYpTBVFapgnnrC4e6ZApihSpG00ilRLOs1cM8eS7hR0f+iwWxU
/rY6huUlXId5mXLUqeDsRcGSCwq6QRaWZMHx/YCfsWBxyse8pqTvVrmwbQfmTsHT02PAluYy4Oqt
1s5YgD7t+h17Ef4n88fvisFDrgMhTW8MF27WEnB+tastiR2fMCBMit2Xz6QVoya5nafCey+dFQpS
xY02HZxTiGA1LaXGuRgnFTsV5RWXHqc73QKzsok9BM3uyJFU9uVxrsL5JJoO16M+jRI775xk9Ky+
HGSmjKraz6lgJtNyM7yOjye+xceN1G7dNnDYCxrWUHzKZVqeh2Mth8fKWQoosporA5LteHLLZJTx
BW2o/89zIqbzHBa4xfM4x8917Npyg4xhLxq+SxcOkGaVT1u9ZHdBN2pypjz+fnA/GG1HC4N8YF7K
GYfiulYq+4uTbeJu4CQuxBx0xJIlT8h491Y7uJ3cTkjwhnXmtFEoE61GgmQ6iiOu0ZusJsB6Xddf
rDzyFMeMKTPVF+oZBCWYHLEmJP5WzYMGppwADbW2EE5dHjG2xG6NhBCN1mReeXJby5XeH8hVbNTV
YvjqfyV4N3Blr25yjse9VftEcREzhrmAdi44hnn4cnohlgHRh5k2ayNmkQMJuhC6EiW978sDSSqt
vh0IAf8xPDxa7TFDiPnTRBK+iv2TOqW8ndm1jrga92SoB7/FqES3kzmMTsUlblplcXuggdoDxEOn
0fWnKhJNp/V69/Ukvum3aAV5DgHRKq18z41qeb0i9rKRo7qIWDP2qbActZuHp+Xa9wgQoYZ0HmwM
M56f3QYgUp11ZTZreHZutIRDUygx2kEB7039tvXI4ZtALuDtjP67dtIK/D5GXf+HZjbF2bNwO8Iy
uCmYkMe8PEEHUgi0GEjEYcV+eSqj66p0b4ylWrDlJU7hN6bk09Ai1auT5lzAfeJGofJuWAeaP7/A
Krspv1uqPd8T4PR/pX1j1htUuf1aBohLDXOqo6G3izl2PTbDIVWwAoYnY4Ic+Rc4b8L056ZioKps
ruLaaX/PXpzXPuac0noGb6soNOKXh5z0CuYQHb1+h+z8J7zkWuO6jil0+Hj/xwwO/3V/rezk8KZz
dLsW5s8Q4rCBx+NsoQ55LnL1PA2gj3CfmbcmNiPYYjCwj63ZH0fo1uQ0xi0WOoJ1YHWBfkPrFgsf
odL07FgpiWmWwflOkA9tmm6uPaFRVeT2w+ZMbtgw8yae7icXw0jnmU3DF87I64iknhoRG0EmpNBP
CJ0toh4cN+o+Sf6mkyZMjfKzKmv1AWJ34E99JCjmWz3916zRxH1GnIpBLdNY0iT7R/rUDx7XQ2bO
72Rkd9Kv8M6qaaGHcH+skdX8d9kxQET6gQFDTJVv5SCNiSd0RRvzRJhEkDn0KtryusfJGdhrmMFq
Ym7SEIAb328c0ROaFWH2KVyVgHPDHqn+N8jpqraBc5ZnuLpkmaPXc/4ygVy03+81On9tCL5vd4gw
SRex9Si1bsmApJzNUmnBh78FdGaeq6zIX6PbIwBdJ0WQcPPdzt89SnUqVO+pXa7l2ddV7shg9iW0
lQDQEzuGPR+w0YfB81Ps8fq0daDFwO59qXB8fjTo7MFWSeJUVxtgEfORuFoPnmOY8BgXrWKNJktL
24VMemA961OUXhVVBDniXRPwG92+CnkOd6ycNkTmIP8k0BSRP9deJBbsDQvHR7E4aKxx3LHnuGNw
LRCf0BMECNM0wpn5qqHBvxYIVnKhROillCD+LTVlL/b26MKvWFlXa1ZBUxL9RS5TxQFjTYa+Qiy5
7uO0+L90C/nxg4vDgQVfe2g9/n/nfEi/1pkTuMjpTTM+F5avG80Pft00n+vUpWNKWmK7xOb8FISp
FMfazE/54e/ZJAFcmdo1BSgFGH7EO5eUOScINZB7T0Coaj9cOJ2ru4n5EqesF5U7NC2qWWRcCWnZ
mpWL599bP4QFdhdvBQgFNMlxgKRWkdBRcUg2H6TSH2b+HSe+wpJ/zz9IMoP+R46uDP9Tdem//hUc
JlubHsPC4RM+mhHQVqfDzFsWRWC0ub2A+9i1Kqsh4BtLrDCHPwuNwmbt3Fm3C2F7EyWkSbYc/1EQ
jkdwz3Wlw4khn1z+pevX8aq3vF1VH3Ys9UxQWUhIb3mzOEDvtwKs0rQGoAE2u/azbFXHfaRULL3J
TamBv7fQCxmFxGrmT0f6pbtE/AzkGY4ZbHTzmyO/fb/B1umoaSfrSF+S9ojEMkZYzFgywhnlPBzo
jUn0elQQf4cvFmAWB35y7dTKeQQUgA88XwEupXLkijPS6B9Eel1gsNn9WSzoetT7pMlxBBxaCQ/h
8cZNCmG2Gu/aXQxt6RhV1SDWXjWKFbBDguYPPjLKxOkX2uFSjZCylqJnKAGXfmRHVYxJ8tLUAtpw
82ByoY6iZrFas3HEmO1PKDuFZEshgjrWFY0C8GGYZZu9Ui0tg9oEhGu92R4hwbhfmoS45XYhU4Pp
4s12TSCmVh+AMx+FfrmcskfMfx5uiau/eK0gT42HU3lrzW4JKYSdlW6sOy4uzj9NZN88XZlOpoOs
//iW8QYS5mVwIOOsXoB1lkhOqimOy6fs0/G1cuFwj+Ip+UZyN7dyLwCPiE4mZrMNMTAJdqOdtOrR
yWLCpaWTAEipfzP19MIlqUh1RcA82BtWtAi/zazvZXGIhzL6bP8RoSu8rUzGnKfPQKmhxMd4fX4R
jyoVOsXD2+XndY+hOeFnKfHl+WMCGzPPO28g/dKmW7yQ5DbUvuP4v2jVNDnNAT+E/tAtKaUL1u7R
8p9UFkbWpVGreNOUz6x7rdmsHn3NvHP3eS4MLtaQqRjnI2CZtAsnp0S8jvrh0wABZq/K8xpeP1Pe
h7fm3qAihp79hbiLdGGwdMBjoqrgDJH9fLZtg7sogOrBWZ8tzEK2VZrdki4J7qfILDvu+QofuS0T
oKjfCo1iA/QDWSGK+PLnGxuiu2EH9nI9+zjPGGvvvyOuqJZ1mTGTD6O6hR2G8JsiuORN3qigBS4P
fElPy19toklOeDI97xPLXcz2h4bBMyfLVE5m0g1X62w3F1P7gABcfaoLTmTbzZMjxKwWIgImX0Em
DT6p/wC2XfF9ODbTFkbOMwTFEIWxp6f8kDDkRbYr/qC8+ksmcqVrSFgj1FDRbXhtxodx/lYGOTS0
rpQmtnFQzX1KpXX1MFGMiz7N+lDS7/zrWleSsz4NF5ET1+uz8eVrSzwWHBI5ZZwX4LroPc/hOkxp
XcGbP1eSyH0jFe5kk85F3V529hz1P3azwSdRkcJkuvZWqbRLN39RCQKy2m3Hz7LPLyR2W750ooNI
Qg0CR+tWDJkd/mGIeeypn/CQzCprv3g2m5M+whi8OOKyrKYuQuDady9CF0x+QbOjkO71QcqM1gj9
p1ehwo8cv5jAXcnkApBhpPGK0lN3I/KmRmTi+KwvHY+ULxNjvnC8o+oXGusCxDhJblMRgb48TVsd
QMoXspIR78aKiqVAHVmapDDSYHS1MKJ+rSeSGR2vZrcBHAup6Y/bUhkezyP4zh0f4BiowcOvVS/f
Jv2m6i0JEV7g2bmdq7af4rxHkR8eqbOd/wymyDUNEtqNqLU/v0w5txGNZyaGY/mT+W1igYAHlpjR
8hVHjRBUzLSSbPbjIEhxoih9mdBl76jwUDSSol1dx3vYDwJExDrKiozCdf2gzyqpo0duHsyrJUzW
k18AZu4GSYzDP32HAfJvkM1kcuNm/QMUYld7Qa9ubcdjuuFyJrTNxbAKj3bW0cJLBk6/FLZsoEk7
7zXNpEPnJRzCPneG3hImhG2GQ6RcoJaqiwpEEHPwTaWy0p2dobtBhRW7xyNVckOdOJYHEhoTZSn9
14Jlxw2RPr8Ni5LEsF0noSEZsw5IuK2BeOHzHdfePcvrWfdpN8aEEx2pLXWrA84AgQ2NH/Rl+hdz
QPgbMfHG3WNFOFzoVhN4mXsSHZ51M6r2p79acFAnq9kyTyc0ccGMBrkDT4RV+y6K7saPIlLLBgF8
EcGf8zfIuOP/ycLSFNxHvTEaGGgR+fnNNTnqvi9cywlwlVyXY36/Y8qYMQKxxPNenlH8CX1kvtOy
ySaFv5il7fwVSfPYDAhhGThMToo/s1mSDYIhSAK0hS/djVUYUeM48PEdB7suJZ+xafcQa7Axx1lz
NrMe6GD1luPBuiAml9xeVX7zrchNghDF1oX0IGC/HpblTNlwfpS9rY+CBKZQ6qzlW9O84esgmz6Y
8wS0qVvSRND9OeEa2ewDi4juMZcwUR1i8FtNXKDtsCB2HfGr3rZRwuQxnwocx6Xx5VFYZ46uNGWh
GxoI/JFkJ/i+rPvciUWKYDHh+uYZ0uyAM+1TXdeySgEKKtnhu3ERCe/YiHrUM1fCHdiyW+pPK8/N
m9nJfzzcZewxXsZ8FE+6Yd83rZZ/AIpPl816w+KoqhCk+A3HTOpGSCXARdeObUwHxenql7hXK9LK
4kIzfBrTw2AgvTKX7GlVrO7R2ba5+72kfljwBKLjIMckZofj3TpxAvO9zKBWWIo2prsvsw7AeD2J
gU0hEnTR8dS43tjB8XkHcXgksVAVxVPHAFemE1GKkjd1x3iMxoPI45QJgXPTbavzlN4eXzBmBVDF
myjlSs1c81l3PRUwXfRTi3zjsMIK8PxDRLNXqkRa+/nZcJ/dOTfv60bcifSTT4eDGsNN9TEPYlxM
43xAAjL0kj/3jz01eojYzQN9ADxVmzFt8AbHdYBRJkaJlyQlbrxEpAeeCl9UKQXDtrKWXP5RHona
krGQr69Xu3KkPxXsLFKC+5KpAWUJvD9dqvQvMW79TA+uICftk2KY22PrG6QjE3ZQfYpCOk6/c+kk
Q8Pifx+H6xyNzInlFdjJIeHKW/8SL2nWtZoWUimcw5vMdkHoF3HOPWlWZoz+Y6Zik3niVZn7rknv
LGFOz6xhZAkXjPuq3mapelamKDkJkmTbh2cUjuR2Niu44ZVZm/fN46/QA5eNJ9sO8CkiljvhYVGv
5aon66daqIJ0Z8L1imA7lK9sEVxhSIDeA1E1DSpxmh+23roqwMboCp8dKKiPCtTTqTw7xTXWATR7
SwjY2k/a0a8s1aQBQSNs5zFqjzqsLifnYFloIrJQ68HU6MOe2ef8E1RWHXyps0izSejPuBOb7AY1
CbUpvlk5ZdjvhpKnXF75U+g/YxWFvjuORVfL7W+FjwkICiHGtquy0bgi55P0vQrsD1ZZxgnMddCH
Do3QrOYwQcu6brRl5XRUE6rRXkjp7R9RkH9r/YhrR9KAtg2rYiLO2T3mHoUSgjzBDMJwHuH4cWFq
RIlKrukxas7wVVC1/d95N068YB75sEuu9L+Za7SQWa/u4aBsRTR9CC0s34mnwL2ef8aNXYQ1132I
JtVfZfT+8nYGguJ8kd2VKk1TbKCaGrMkwulInZm3Zsazh3qDP7S/zFcoD3lNIIVIq5O4HVbLth3n
sTnlXj+x4/RrwoR4kU8t8i563O+fnMxjH8E4F6z+LBSHFX+oc8eO5u2ego+FxXUqxuJwa58QojwG
rDhEOznft9kkNbYVAydToHbmnZJKHmoiPBeeUCn7kDAscbC/chFwiRmZtCDHA/1ugAnYgZS0ZMsL
YkTMrAwdw/8nqdmtfMHaHUPaq1J7EhWpC6U1ZUcUvOHnqIKZGjN3WeS1/YHNsgIxZvHadY6hGpE5
yyd3RLCAEeJ/6aodWP7SHuYYTcbusmJ/NYTeOeaZZxwRVB+NL1cBOsWjo08I+vf6qmc94EKnGHD1
EZgconofCBAf/+5+8faYIO7gcstoWAt8ZobY/wKqIb0P1ubzTedd4VykeEDJvuXkEtGOziiaw1ov
Tdq+6I/o/gn7aGq8+F8pvE2v4PG6ea47Dz7Q1EgMFO7hBFSlkgqylEvN0n6dwwV8J28YpbHpdjy2
W3o9T2SVBupKKqTUBvsU21XlRimuMUPslMO/OH44hFf85xvfYqM9cd2AqYBIvTQG0rs4ZT40iJ4r
Ht8cow/sJ3yIQ7HnGBia0VO16ZvhH4NQ7mJizB61EiThzupPbL855Mzkd9r087TIHQBTrLMK/JMF
8lyI75QYIel5NHprnsL0IPsrMfNrfAM96tXF4i/IRRVCQ17lcBqE1XwRPdV2vUtSWyB1qdFVTTz6
6Lzhphw2L7d/73TZwsCdaULN4NfG0G74EWOBwiTUUo9MwCRaHqIr3ujA7urXV+Aai3uKqeV46XvV
cz3EMyIDBf6EbahlNL3aNYeHcsQRXsMais1P4BaXAn9odT/2ZkguDH6gy2vbZECAaebe1dhho7fy
j5owP7CDoki2L4G5/SPUJOKPF+pSOCBkvVddHvdBVmzhuCzTo+16p0xU1m6JvqmghohcHOZ62R5o
accIFKBnyZdjfk37rAXIF/MK061YbH03VCUhw+5LBUop2SW+/BCR6rBElakS98uKugOvoO2fsZgv
TTQoFKvNp2YQ3cSoeaVwDSskeAKPKZeXCM6trNIu35FlfIN4Qdk4f0hqno9T+v6Jg3fUhXUZ2Lsc
VijqUdf1BWEuHJ+ne9OXpLwh4F8YK3+ZkDyb1dC67HkqUXju5Vlx0p+Ge55PQjlpnpk6Y3CtgR2l
0x6Ds5Anu9wrnxqMOifN0SshO1/3sn2VswNWnoGeyaoDFU6l9THSfA22FA1etpLR9Mt1VrHfxPEj
SN3+7iiOELRJXzWzKgjyEjVxlF0BkTjSou2wJE33zaN7EP1M7GgJrmc4+9nWufnxuS8JHatv0MCx
bxruF4al5Cylyn8TbXb/7ZDMizzuAperJL3nlFTHtkwqxBJIvrfRk9Onr51LHzGkxNqDUoEPUsTf
gOB7K4ZOkrrPUVXWcfnmybEEglSjnOpC09QGefmghlh4ewNaRMU0GCmW+cGbDgQNhvWBnQvxyO5s
Nk6EUc+gVV/wFR/1ITqSLhspRruN3WXF5EQ8SEhtw+VMuhtYeXEnTf5YrUOiMWpFMVmprP+PuBow
C8ZZdO2Ywid2L3VILvFhJ2vNYxOh1xTM64SzZU3pfNTQ5vJk0T4OQ03Phz7hy2l7bQAlss3FUupH
7pUPqn7ybrNkpufguoQWI8mCONcXcWQJjkYFxlw4cJRhqwDiqTc0CsoQ+Tho2xmzYRYb/b1HRRrh
CH/cxgfRritAftQap+KymMW9AzUeRfGf8GbQW/VWyGG6mfDL/9s9sHoqXOeiC6wNhoVeC5I/hfMr
/b9sQodfUTQ2dSt0IL7nnyzjQ8fqH/gdz1s7abvOhrbaKB0D3x0/bVKu9sZCTDU+Hg8RZR2MGKPY
Th4PNn2mfsSN1eGWxytgc304pLmv3ZT5wyYnwzMTx9NNXaZheqIlt5E+kyDYIG+iKeTa6jryi1F9
CjhPRyHOfeVjIGxYSHqvYdvkr7/lHVKe+urbIttpmoLPoX/ERBkHEsslDQjA90veNGdLmf/sTAuk
cUFVZouAGKZw30FNMsybbez+y5CsD5nvYT3SIZvjhIz0BTbKVM3nZlEwjr2ooHJTL+Lmek6sQMpa
+8C+xkfkWxLxc/mzcJevuIMWxKqUTlxwggJjrF3WD7FCE4uh2lhqEletFvYOvn58szx4l3kRb5Io
DpyDmgF/S7cbR8A2SevzT1FBQWbu3eoCVelLqeHrAWTaNoOjHFuIjCCQDkIg+DLj//9anXwlKQeG
FxzbL8FruWxJeFSg0M4RTeZXXoMOTUXEExdSV8MUZ1HHHRFDCCy8HdkXLp9gXh/+XbCqM/bvQ/cj
fZjCq7awxRH5i5weweeqd9kCX0CEiFPmu+zy9FSsXg04jDdX3htq2Q8KXJ2R5UljEJANVT7vb1ia
YSrSfrpiIjpKWiR74T/Hr/nF9eHT6J7dUz9/jpe7aG6o14Vvp0M1VPDpc3ywqwzYkbqgEYQ7JmxO
L9HkbyTRCGOCgomFiBMwqQ8XRLq6Fw4xkfkvw/a/dtIHSGzfNTXt82gb7I5w5dztIBkj64zNJwTL
MtEM60o+Wpy7K9cHHov6/ZuMizNoPHSqMAxc3kBBZQVc6sVkWkKQVU2Pi21HKuYgUFB0g+w8v3QQ
/M2gbnmsrc4swkkrzW9hJWYLG3/1KVX8NAQ2IOqdIRbCgNLmLg/3VACx/itUonzbCGawiPPT8yIJ
ST7ff4+/SQmNvhSE9QDQzJ8E0xYp5QXD8DEKaB06K7IELUog3t+BpsZ0tHFWvbabCg4LMS/EA5dC
IIGumQgwyG+kw0bjBPkEP3v70xFqogOdHecfjhnku+MtAhWorvEfYHg3RWcEFbqQXMsDj/XWH6le
UOAwScyQLkKd6hJH2R0d1aGBoyb2N9wP8IMcCVgKmsEgW/orev9PT8NcQv9NP8N3uw1HtQob2hsw
BhzH7btCqFwgbYnTlaTIbS7QkvY7IBuTMTf+n8nMsEqKpavrCjMreq53sj8ucSTLKHHqgZmubmEO
+G0KSrDHGS223LlRAkZF1QSfzAvqSa5amycyTIG+uIJ38Y6dYNqW9HAppJF9M2Ak7MwOoDkYo2m/
WKU9RMOX45FjfriwkdlhYeKYQLMnZe5YzVXJ+Ho2cnD15397Ldi162kbYSE9wlzoR0y5px+Pt6lT
QtWrGIaFOrKn9FYQ3379iXOPJSx4N0cT4ER3EPI2HOHpSCiXHzFQAQuRcHVDq15v1Hhw3yaW3CDe
AJIPVcrGtJHwVp9Lfoal32nfI8hs4XZdG3VBBBi+/DVC9+IAbYYMjm7mnSmcVawfPDauxBctZDEZ
g3B9At0nKT4v7fKeOpUa6njFhGEcPM8n0YJCIGVq9DbDzIR3X/b/xlSQSCfNZYFkiaAfPiPgmhnj
zvcmckhkNF6YQMjJwZgTBr5cOeJ+ctXgryusiN4CZmgStCY521mMQ+/p2dEbGjvByOBxNpWqvT65
i+movjw8SDwlZiml8D/hnU3vqYELebQqqwyj3B6V5r6UDO/BKxUHtzxsnxLCENYWgguYU423o9ca
SQ7CxxxoG++/Callh4eB/ZJRsAcAevBu+zjSmGdAD1Q6ZqCzvGDZJRaC20htNgK11zhoKkSpFbmq
g9Qezxzv3qEcAIe1aKaIAgdR8U6wk8LJbUVG6KsniSKBNccR7uG6BvyfA59MkTYX485UCx9cb9P8
t1mVw3kzvOeFrOGXLhQbH2PMD9XV+Q2x9+NrpFfLbTgCR9Kl+QS2I/xPwVnPqyJTb7lshC7LRBTX
3pAbB8J3Bm4qed6S++XoJZbjtdD/jy8LglvADgupF6V6g27T+eYjlLHrsPhihX62iA1rY/qUtF+2
Xo2zbxgF+CybqolPldUAxh6NSj9HaJaCHTUu4x9wLtGDMrQmGmPbR0cR+CqoeFei8oEttCUTjMoq
gq5kR4vwk6XAuGmd8kuPbKP6nxWOfht8d3+/+GGolWqFfxN406jx8BOAmgC8aMupK3ejIHYLBjYB
XlKAvVte/Z0hMrXeHnh0rIQsACpGMmioMEyL4lDHT1sNEZeSEQTxJlmqzA3aSfN1+b07ISNIR/se
HlYPbvVeOLQFU0I8xW12FyOb5BiPwozFTlAXJXUt9ii12dXIR75D13VLg74PcJj7yeFANWv2E1P4
lDK8Z7/N2DB7lA/zPx1v/EsI2t7WiaUy95H11TbDb9ZuHwYnkGacVa07iI9kMaSyiFoVxF7BnC8r
VOj3vzRWMNcI7/j3Ms49jD23RECWI4cvyPzD2fzbOUt5taBe0LPeGYvbBK0eTc4aC5/nqjFB6t2L
tbtRYkbnMmbR3bX6uwcRKMoPaiI/E9l2aYhEE6IMtbOx0qY9jLFKchHDJevxNsNPwP+gI7dMxN76
GhVjNrff8S40exsbtUUaFSe+9v04L9cPcPbS3gClSiRqRvGniqp68z3LGU8O3CMs67SicITVtvPZ
mHjkpFcSzbqvtjEN72p86vKmOjCQzaIELUeon38ik/ZHSFshWsXJOKtDUdOBAQZdHG832W7QqikS
1oeRPAhCI1mfyAoKXKDfFXpkBlxjAPJzJeEbziotGw32YGe+lKd6MLVjxWW9t3H1IFtghHnijsoN
TWgpAwhfbmhcvsDevGLUeHIqgFjeDut24LL3eJ30D2uZrzM7NhJ+MJ0hpih4/AkN2tUBGp2NhsKp
STK/xKUWXVNH7quWhZc1dYW3gtTVZbpijYQSW8rTiSbJxMnbHk6G/gykIrkc2XBPbAIJDjMoLJvx
Rv3DNWpP3nn0jI1EecSo7TyhG9NW1WPDlReJceItrjryJAX0kCGUR8vF2QhxLqcUDPZVSSE0SH2O
jykutNE/sorEafPu/EiTxc6IK/2b3UWwzn0zwh9aZ910IltiVk0tJt7DqHCSt2Q8pXbzu9/I3Hql
7AeCgfB9HL2RqzdRCwqsCXedgs8XgwxmVuIu1aPwFxHifsGvzIc6atSvaXBxPnrT5ISneDRbftK+
h6aWqSf29DZ8RG8HrkrlID38+VTVFxrF1KSo1jw9R1d9dKNbUPtm96msKYFBkoX9PXZX8rZHYVxX
+rc5+ae/h9eyoX/obnZNlS7XIg9uOwQ/Sz71GtXuA6x01vnr3fRwC3QAzlJi8M/mAxyWE1DybAg3
O/S5Ys9kilB9L1CFq8h/UjmAaTidi07gb730IpzvBEjPy9RfUl1qOxNnkVOaonWZgi/KAYoNe70S
dUpXPxlncyrlVRnCkEpn6TTl96yfu/nkUQtWJejsq0mv9CxhRu2llawv8hf/kKBsk1Fwl75W2f7/
dYZAXChdtkKlJEnQKNGN33iR1G9NRy9uDUx/HE6ZaMT0oeC9E5n9uiIJbWHfOmQDUlXL+RP+UqR2
BJu9guIIYpxCiRZtTfuj7IfMRKJ4f2BtZnN0H+wMvLxiE09zjWbS7fiRpfpdfa7RJI6krC4xCOAM
NfxnX7Hmy05QuuVuwZt+f4HW4orkEwrtio+BNYD6aKzHzZoS+o83cmXUC6WtMyHyZoPwisFEpthB
TttgNjfx88Hg1K/bp34eQoocRKOdxH0pok8sJy3dSCqFwcpcsvnnDcp+ntOWaE9/8BNqLDNWnfcU
EkZ2IHQ6sW5ZxzOoC7dVL/OfBvM84mm10gq8bmapPOvo6rTbEAXHCHxQjr72dIKxitdJM8fJK6i3
uCq8qiea3ievFrSa48KTgtw93UMKPmev33bBedcNThd9dq8Jwu4vfuPG+tBu0qx3SIku2SwNiTDq
C0RE+bVRdgz4IzLAcVITm6BGV0LqDowjJhUaLFjMQj40EP1Qphq8NTnAv0lad+LxlLKS/2Lr/kCJ
VsKVa3SBUdYRm/JfU4Obwl3bQTSw/W/pfKb/tiNFPw1O4RmynQINaGTCWVUimOoe+zwulBE0F8Pt
oEqrKr/LI5Rn/wbHlLug9ERGIESUpxQUdxNl0oER4MQSKB8CLQEqFYfrFJZmpDiNog2TTwNIQ3XC
AhCSLlfzpu5ORiu8OfFT9m7RBvs82kwp7PUWc/gKW93eCPBINoIXaJ553bDZyBBM8o/yQa88ai5w
dKsHfeggZNVtHCmdv9CQMEFpriedN3y/XG8kRkx44pel9RryHnClTr+vsa4d0Btqg0GNpyi/+xbE
Rr0OHDlPpAbo6zry2LuiqKhHPIz7NqrIHaOOjrtRoRjPeIJ34kHfP6OrTnbhRKisEYS1Gfii6BxI
+y6KLo5s7dTZ6Be2/j9xUd1Dvaf6oJMm3ffPX6G5zHhKMFpcQOrMtjt0SOTBkYvcS5UHvnfk8NHr
5ZUGBGhABlU/oTpCRsIjdZaWVyeQsmmHGGi4ZqBPQIg/hEgzN31MES203WabHkbYpwg8PrDkIqWX
Sb+9rvKmC5jzzHcNkMqPfg5tFrSf1ArU04qUBNf3SpypRHTX5y36TIUoCRNL+zqW7c3MwofnShim
mO7WJXvFno2LyNuGZagTwI/MAXAGmUvN3YIi00+2cqFEfLjkZLwrGO6Kqv84AUTp4dr7g7F6iif3
aN0h4P/eE6yHDf3Svz2DSnpU+lhFnNBFg0S7W3glQvRPkh8xMZAYEiRhp0SWlrTR9WZkmXAi09Ws
Q4pbUS2MHTCjfmIjqTF5n6G/n7lBuytS/06CzkBgtvrF9cAxxz439DXVWSN6uX5y2cMsWg4MCtYU
iVQbYGNnYjGwFromerZgLNtmwnc6mJFIs1VaU3ntMZiOGN/N4Nl3D03/SYSZS2gv6T2reJBojQM7
Klyzgnj0/gj+yM05MxC8v9cZ0M8cNzr5ZC0df3ipQlDUBbfBbSp9fogDXR2Lj2LbAcJEgFug2GXc
RejhOz7BtqdeyTjEkXMrt3FEdC8TzPcMlaO7diuGhoILN7KAMXlsHJwpQqcHyQTImnAPwXupPiQ7
0lsf1+y4UiTUNbeupKvMPQiebvd1y9ao79IR5CCkgztwKabw/ylnqyL12nyiUJfCANY8Iq4SZqTK
fDcbE4RL4wmHnmEU00qtc0ktXBB3RuwrskT8eGJOLbU6Ob0pEXSxR9EZNOJah/Jeo+IjOdpYW54Y
nONKIXOAe2P0n1aWI+6hqxaVpGIe/kvCtgo66KmV+UuPeScQPZeWkbWmf3tot/+w+kTssJVd7XD5
piQ+uMwbsmsTg3/5U/7v4/c511t6q6eo+uF8Q+KDHpJNnTW6IcsjwhvixWiM8EhCcaaEGsFwNxQt
Lktarnlqbde1fZN6Ane5T2uWM4YGLDBrmrZEpl7dUw9G18DB+U6cTDpFihjIUUTgHhoxV2FHNdLN
e+xKRQ10k8YG7vWbmUSVFZTFnHtgo7AS+bLi3kDOwuqM9KJKfb1GtHM7hU6FdRMlVWj/0zL9MY81
K4hFGdQOh3A7u1CvNO4kmAvfChHT2aZvqowKxYuQnEa3z4EbEyynd4i0ICJHaG9tZnFpGeJm+Y0C
0kPb+LgwHBkdVuz7qLIs4/Of83FHzK15ofUUHM7Vz4pCJfztdNRtoED+exocgrXqiyzHBp+VweGt
Z9jLOkGr9JBqjlnSM326C5Zzyaro+yNe7izn/F+BEpVhdO8wQhkakc1GRHteTPFtJQTwxfI59G7e
AEs+hOFu/nrN0Bwd9UJn4eOkq9tTg8r3qIrBm3AoRMPeCASK0jSn37zdlv/i6tRr3JIPYN10h+YC
ZrTTato3Az3YSXTRYP9uueP0e0NFru6I9+wqLoc2tsRFnVUmlo1GZMBIs1Z2ix6t5svvoRlRNkHJ
cXvfmO205Qoz5a+Z2dPGQo7XOW5YfobHirbc/Bn3fLZLMRUMFxXxbArFRqVPdPGLVJmmhoaSg/gg
4Irm4uVD7ebasUTi/v6oY4mIIM5se5iFWomfRvWXUiAC7H/oQvKdtA79xhYfPv6bUtsAmcYj2IT9
Kth+3rJlxiRMcdVVmObsLgWHzlobg5cX8R4TXWUjLt+EPwSmHakl/jjYte5birvRVu8uvYt33IzH
WJK9nKa+yUpw7kRPCYCiuz7HtE5+62btqoxtZd6QPiMeN8O1Xrh8cEIjwrRqU00J0Aq0Ot3PkmcK
W7/9vIsW4Pz5Hg3uL1hBs8lBQ2oslnDOWJmBANvgq1xRwO5iqDHSw9+ydesQMBTy8iI2HLye/Ud8
g5/fTZFHDvLCURbMRHWGbMrvYKKjus78cjRV4ZFPQ/7AxkMquAtBEZbJZuD1Ozw6+8rR7BkdYVIC
gU4VL/zhkYknXYkdm++sQQbzWbd5ynehL/ONwvr5hLIZI2muWjpVb8lbryVBwXbJhIFkV6cOzUlK
xzM1JqQrUsJWDhKaxndsDl76KToQiQQz79okN7CFMtOj908T8lix2M6I7wP9XRLWArVxVHomFrga
JnD5F0ArX5batQrLmP6loBdHfjIzvk8dbrr4LpN7DgRj/54grHQ/i8UgbMZXsvA39n2KdnLaHFue
FzWOo3ISNOIAadc4n6lv1cR4BE37RD9hfJHanpsqlgzI8SYovIhOD8TOxFSsqOQpdtM7ikUFuaZW
ripyhAQiKdC8YfOno4E5dvUmAdXDG8wkUyue2j8CDLlqqmZWceOhG2FXXycvvilNqCd//XySmTPn
745CzUKNYMYAFBLIByTGpyI1UruyqvAUjqW54EyrPgB4m+TKtdY7tnubfiPDaR7/d7DpwacWvyCH
cYnNmNVtJHPxti3773uOrpyKikiOksd1CalKhtvz4jU9H/tfzW3gO8SMHAAWmrggYXVB1K9qeLdl
9yyTHk4vBD4rn5cFodKYQCnOOd1s5hPZRZgu7ZSZOgAK6FmgsEQ4FlgKioFkxWnvobCmc8pRZfbK
B13nUAuQ8QWvTtWRgwU2BHvJrRpakrs5NREEkvoso9WwrRYqo7R4nBkoEsWcL7CFkHCWCzw8AtX9
r3eEmLeb7CqhQ3Y8TTjnnHJIh/8E98zukuzXl1X3cS+H4XmPSIMBFrTUmlaocB32B3FH5n072gh5
6H9v/+DGjTh0EMukZOi/mEndevOavs7q13HoJT4lgoKyyW8/DF97rq/iKRcz8SIedLg0ydxR9sxZ
y+nLSzgJqXeMs49cTG67EHqy23H43AQTZdxwYJg+y3FHkqBx/FTzSW73vk4fxPJKqPVMwunmbRW2
hwmu+saUrpk3AzpTcgyTBw5WPcE3E/HSL4Li6Nc8CZpjOZA5WDZFQZC9o/CkydeLIAOqV79vM1pg
kCG73RAHRtnPfAcHOmReicw0NNuZ21uvOiYen5woEgkbpk5PoePaDcOE2uexVCaazWgc0sqSiiJ2
JfOu7C36vAUoLQc4lmtqOadwcAWg1pmKhWuORJ1tq+8/OVNwUbVDeZyiUjgiqT7yaM3TqDh0AOZ3
L5MXEHFBs1LdmW6xQg+2nRFLMcExQ+RSikEERBgCNMmtBMxLUe1AlNVYECBvVOVV9j/YbulAWaSB
fL2V+ZosqctyFqSDtELnlLgEhmj+BzfStfX2mjTp9lw3OMfuAhMQdCLz61mDXFlT3B71TeSHuaHy
4p3a1So6n1XSGzi7ZaPN3u2lvdAZO7bwxMchC3rcDlyiVTaaYQcztzCORMdXvre9yhog5ed/T5Lg
v8pGtR39EDomyO/VLDSUmdIDtjYiXRVWEjEpYlF6jF0Z49YYnK8wh8EAaDF4QlmbhB4hLbVfAvKn
4h3RO2K1cohg5cdsrIuDa++jpmKMc8P/HcghY6pJpYNd68yfZ71m2qsk/GfitmmDxkTYqXPM3dAF
lo9sAxmrFDANAS/PkP1HQgS1jFHql9E+y1YWtInpYdIKHsK4ovvkmLBne3zxzVaYCFdgxQCFk2yZ
UNBWT+MwfkrXh0+0SIOvfNkKCoU/mXXrxOW/hwpBI7E+p44DvxGS7TM4swG448EjXuIuhicWhfnl
n0MfPsUZv41UZ3gNfyYA7GoRYChXhF3qRxeZhrx/DOFVNz9tG2NA7woo16ZDbhLagUfqaLKrU7jn
uY7nVUxErOhphEI+7dNgTM2Ejv8IWV9LDxA3msekolup8XKMcMsYwrkp8IIiR7XClg7fQejrsILl
Nw4GBgqS34qHKZ7q9mUYgGyNGNcedB7seWZjobozUYQuC9zpbQMQE+DwuBayDu56e3itgeuRdNLx
A2P+p//3KXCVahtRfVQ6a4mXPvFobOaMjtuIX2y763XYv/dNUQXJvU9ynMIaLFYoZNZKm2FvBaeP
cG4x4qnOnIieJ1ZanYZHqXOCkLu5SJctIDaEKD15su9AoCBPXHgRLkga2Hq6svIu9OPWgyHf5/fB
jUlOWtB+baeNb3PkC/9fz0djsp7OpO/TWmxOnO0HDXB9viAAtZ9BOxRZbjGNCgH/xoB0qF6WC3zW
Um7NvYIzmm97f+YCaesMywR2EcdSWqa5E+sSB9WSUYSHmOXI/407UHFRelg9SiT+zSphHjyPBd+5
VIWCBkTBHB3z9pKEd5qtDG2h8vQkaYnaqMZ0gYG42c3EQUQF/y6st0nEboJuYfYUHytvSwmhnRMv
gJnJg7KIt4QisasPTKW2Ca2JZmYiCz3plIvPO9y35Vdqc+pwk+hX+x6w1kKXSQzrdLpKQgDfvZov
QUPSGlDHEjd+dZsek9rXRRinQfE/b9p5thStQL31KyXuKZsCfDeXYjh91Nebg1GCQnvVE4iKBq/Y
JwWpzPhayno3Z2t+rv+PxNK78ZX1pVinhYl0lE+QudsNOlK6gZqIM1McvRK1feFtzeasgZ2MKeXI
z1IWcv0MQ+Gj5obekM6Ayc96jEsDNK7wcNTRvN1pkAVNY8J4YJoM1OIXYPv573xcceA7vNCjT4Qh
As9vY+4P20j+EcZEMv5oXjCB+JZsMJJvF1qfpmvryxKflbe8MeopG8uJXVaeVaO2kCfVTRMqusva
LSt9BgWpxJAgIQn3JUihdTUCG00LlQavI8dfz002lxIU+3MTXY9HDpdfQ0COBD81b0U+vTruSdZG
TwpPlGEdEE+Ipx8PkmdXo748A+RoDspcRFMAjIZMAO/En4LtStXGj3v6OUqwvVqWRGPt7bO1owwM
9eM3Vd/r8mtHIbGZkmOAKCqD8LDIs3bQZgn8bypzZRXf0V3DgVvwN89hZ820K3KcU1JXXcjNeUe/
xfZBpiTiIg2wGnKqYSKAbXAvhpsByxxOXprWFnch1HLtsTDts1OtJNH5sahqAOgQCM0YInYmmLKm
i238amfN3DRNzu2dHkXqkFTvKSWVZNOEK+dYffT4/kGk4bP6QPlFTRYfGxeRds7w3tVsGob2XXBC
RdILSJRwXGYH7k0KvvcMgN3GetSRllcd0cQB1NN2jEe7OP//BOSFoNX7GnrNhNuDtkMKjewYJpqn
FaNCxmojw53rYY/hUgHlrlyMa+8hHLS2Bn6AnBw4XwrzUKfUqGC15T8uJAdK372izmDO4DdZLlmZ
PIfEuhWWbgaKasFpyHmcXMUfP3p6wC51FTgqxcQrRSktavIxhcJNWX366KzgvO27kxzyShqBz+ss
LVZGm6BFmKGZetTpWssSjRQsvaDAom2ENKOICU7putic2ebPwLkzFj6wNQ3XApR3VMQWx0p+p0xV
iFGCE2p+q4uVzzk1gRFZ5Ajxi+a1ZVte42N++ljlBZ7beh7mHCYlEq+9Mr3c6Q1y79qW8EOgBgvJ
j1QYqgSfCWbj8biMmRl6eyMMqiP1mKszU1wqKNy+MgoBkrcWiVCneJFDIRPSRVTXETeS+e0oWwvL
sykNrJ0vtkcsdMX4WBIhsxzrG0dR0P3DTTmhvD/CWsvUEEK+lZnAyslL8JcbeBqBn76dYqjxQDSv
j3INUry0lW7yQRXqIihIDKYW9oAZQzt69pB0TCmfkGx/MbsDxuHGVrsOw3f4pWv4gjZ7YF/c/lzi
u1nx06MDGiWc7C04VHWlUF3u41Q4sFFn2SwQMG+7YERL02fLg6124khEdKnjrvz+DhMC9GMf1M1M
WS4MLUNPzJKhhXDyswxWinIpS/VmCAsLhJLisbNQnu+6rgVzxNOU3O8c5Tc9ay5UK0vHXO01MDCn
MhEYDw0E6PweE9GgisMsQRWM4wQ685ijat8QRdvBXJ+KBvdW0Dgz6BB/QnMRYVYZOgNXwtd/mb53
5NNYXCWkLDWpHvdyYXlIakVQth/fCjkoAuPPRcftTBUctN3HUJKMVJTj+5nFSB6mQCLhSONHxtET
3WPjVucMuimS6kCNOzGzHZTFDcAieaRzHu1rWI4wYEUZnLWXs+ekf93WAXQaWT/TFYhs4nvPt2a3
flU2samF758rTvG6x16TEVMFexyIHp33aQWbf3OoIrUCF7IP3su0e61QoaDx8f2nlxaQ51hGo1sg
h5de4YLdgPSbpQx7yqlU1tot+HUWfiV1u/x/bTz+DdyMRaRm9xu/Wm5oCZtkrC72iB4n+01EVnh6
UHS7L4b5zy248KD0p1spoiI7LhQ5R2gXf5teoArxG05X+QHy1j35UtW5cgP8E4CDfaDF1Ih5R8dW
u6P3trKj9IKXQExMqNlsd4amjzW4WpQtnXCbERUhtG1kd5NVlNm1n5UEijGoCCTQC2G5GuOU3mZU
5bsHTX1S3YLJjEw7zjhz4tUELBpawF5bXmzTk+rr6btUk0a3P1mwvG9BgiHm3CR2eRZEViBEfEqM
ASfcaOQlFYpeMPj3BJGFuhLCepmsN34jYxZwusuq+gevjsSQprlFSYeWqv7RxzC1w6yc+OpiE3mH
MXPgbBuZXTIu+d988rwpeoZnZxvQwrHwrvrwQoo7jd+u/G14dQ68S7y5VqBymgtRJAFwNIXqcjP6
BKy2irdc2FUOx1tnf5OG0xU6yAjonjicONfCZy1woK4VINoxwkfcIDtdah3pi2p7ekNiVI+RL5Vu
uJeLn6b3kUqnCGSLETJgCx4GKhDSEEIzdSPXktsvCWBrF7t+7h81V7xqgmvVPpjpdLrl7Zt72igg
G/dMQ7B02b5Gwr8n/5Uw9CfeuQcOjOhZDl+KwNvtvZYodcQYj/m61b9DlC29EWQjblEbKQbIomGz
NTgEkepkvIwaNwcAcqCNFegwnK/VBfXBVdXTq7MVi0vHmcZw06ZsqdAbo3XYCp8pO9uL5jDzKUft
JIK+MJnJ8EXKOfVuf6d4yJtKcyrmtkOZMi5OE0HmUhNXU+iEp0SCB0eyuWxotH1vSjjBtEOPTvec
TK2akyWE51F6WiO/GZ78HkFvP/OcwtEnFP8d83kxjIqixgR5ODb2Ex55k1rAM5yq1COF5IzLyoK5
uylexr5B4EgRIUfu1cFA2bjyGH71GOE5Kni826c6juQ54ApS0l5/x+nCWUlxpeShH1LDzn39szpG
0VYAcJitStFSUAwwzQz5JJdPq70UJt/Dk14lpFykeeMtx/fupjOYtL6O5hlC/3mbOpP8/8npT6tQ
Wwt/zFx8UlPKiqOGZWduCFV+mDf54M7X1ULz6od/rBE+6aAnETiJVyz4rDeUZu0rEhkACQ0iii0K
QsONeu78dbPMwXm9xUy0oV9YGiCeT2RqYZ5bYrD9N4RopmCzvL+CGJHXDU8DDxqc3nSIthQlRa3J
bYkRQT+kfA6d/PyRSU2lXfOqjoT6YRcM5rqTK07obkS354rOebNl5kJoXfh8GL39ot6UgaRsJdAz
R+r4m0dhNRZHo3plogEmYl/DnZO7tuR/mwAbKgPvNPMqoE0QgJwYjrq0llJK3A+o13Jf70CToO9J
QbINVFsyaL2XSmV7P2bkzvtOtG88etnRehiRchYcXSOQu2i4g5oZPl3GQpMRFbU+OB6kWuMYw6C+
sMNVYtXyv8lLViA9UqoTiV6Ewyo1ic1o20XvR2qy13t/Mtp6LA69eQm3AXgyZweXDkGYwfuGAwZF
vllaoVD9KCLTyBuzHEeB3Rk0PGI2tZ03txsoL5iiBw7Y0I98L1ab0hfw2Q7JHDC/7lfJQPe5oxBv
M8TSB4m9JdLlqnR/vQtlp5do1rOsxZe0CsiqrCWCz3WSL4O0AaQxabRyD1ycm/NV9UyXONjzGcfL
IyNXUTiW3BV48V5L09tq7WTnFsNNR7oOSkrCw4RoUMzF1lL5TkOke8JaEDy8TKEJS0x45Kd/RIEw
0uAMwjwZqCEVtqS01c+/tUcrAQxeL6V75W8ZJ6CvhO0t0Lxo1IarmklYrdZPsuKaBlvC+vTheig0
WY7gN5hD3JxCamKADWfvfFSrSWG8RV2acpMI21KuiJ8tXqYMI9bRuB+9pUI9ZWZldi69L+tEAWGL
tvWO+0opKsDGtBHqUYSy8364GEZ6p6SNXcXjC6LSs9QSDuM2k1R4mkTXqnQqyk7J46ymgHPpFF5A
lRHD2+JDgQ9BUsEhW8Q9otJug/i8jXITpmaupqPCRN7I/8Os3DcYUTKo409GHSAIUPUJ5zVudfUL
9QeB6tA8iKwo7Ux7OXRsM/rRP6qkDmyda1SoXxUVZ1xyl/2nKscYtXldVzBWydY+vd3CLtOS0wKk
CI+zxB/JnLJyCyqpu1C1cdvjAWRp/1+D+SvrhOHt2QHsCgTRNfXvP54fj4zJBxyF2DfiReIb4OXv
+/4wnCCXNQzBvw580WIWAnyfk3XASG4fKrGKlLVKDYYm6ci/WMZevYu+vmq3m55S5JZUKnzGwxDO
2bpVU5J/fbN4k2CEKN1Urk7WP8SdhS9lr8XU/73ovJ4XG4eH1BAM5OCYIvLygLGFgLVnIAKVgD8f
oJK5k/Uk6veacDFTgGjJ6wa+Xg81JpcQbQ8Lk7WLgIrsihckFxeRY0o7mEtvVmIAmgQpqvj2dgOW
BOMMw0ZUYFwP7MdmwAM1ETMzeAPOWQEcI19kzxRerwRbuZj/w6dQ2yAd7Zy6CNkhteMFcHbuT7dd
SlhCaK3oJFqW6tGsJr9aL1SBRo1hry9IIisXE+0wfkesPtKSgTLstQVooVX8ZjMgEnyZ2wwyq/mt
nEUC3z5mV3lRgvUVcWvHXlTuOY8bVLcQTMymStG5bsad53SlmKdl3YpwaWVIjPFjCDKaaF3wC0WE
XowXtshpOo0VajcRlrH5njheu6M1C2dTdEGv4dFyCwb8sSf2RhqOtHHuYgh0nu7bsZCVf2FIaINb
STeOd5jCwFthT+RysfElxalfmXzmoCrVWpd0IdJFBr57gDJHF6LSa6PlXNnHk5/j7GzlL1eg9Lw5
p0vQX05KIDjkUwdtPiGBUnaYbwuuY+RBP8WgwHLhH7U71DGUdqtigT2ZadBbOfmSQSbcsHH9WJf6
f/+FjFCoYJiOWD1c35hWnKFyLpGATk+6yhA8tbM+F8xkSNp8/++2TLelNZd381Zdh+xb/7Mw3vhY
+MtxFc3qYgFRRcxRXqE5QO/kJQE3DAZ2/ywsk/GTMqGUkGer4YOIOn30FknmAtV7oZF86Ijmvuzg
OiDd5mb8wY7vuVtoqD+3xMhnnr2uD4/m/78IiJlbTUuQXpgDSaioQKj8oFo8AAmXT46oJf1IWe6N
pqW7N7mi3Q/KbsbIFsWswms9gDEovwtdkOacZ2lkgRJ1quBjPm6Uf3ni1PzvFLi+fR2+/UdFNisv
zZCJ4MA1EuCWq9v2KBml6fzgZi6nKDChTa9wRk0SgFBU2lolYFz1gwx8b6uJhgPe1OkvDRxoSNz1
870sXw3aCBX8VMiQu1of/X8aniggN2Ca4bEH2+OMT2JX8AFbogRnja7749mC0sMEWttng1ptJZOr
hjTYUxHjFbJvRM55P+p/aKO/eW9nv7c3lgwu8wb8IGRkgzbjH5inKtE5qFkqNsRRK6mJ2F2/GR/E
Gvha3fOVt7jInVX5mPiwE3hNQ1R1MeOxtzufY5yW1dl2kTaZ0BEi6HZ80jvUJmcHAo6JDWbKeN1S
Rx4AxW/zpAQBxzeMaMiX3cfzpY3FYnJRsoXXUd68Dm0FrUY516ptw4hCNuKe9u0RyMjE83+g1h/D
dBzuHZKmTfDg92ltcWRYjLae7+tQUhx5f5qH1zY+RAqEr2AVq/l2nSdigkKURQ16mPsRsbBMr7p4
57V7BawdKAjZCXEcKlLKgSgVhMQ4P8qllHuW78X9vjQhjchWxjJ481TI2uRi0YNX9u7RLGITd0yS
FpDI7195kIOxdzWDWkflMOrGPu+mvIEPrF9kSSxeg8kCPXxjlKVu6il+tEIvF1nkVoCjci5WhMxC
yeDqWpA0kGoNO4QLmF5Sqx2+hvUbTG9i3xIJHEXxVrd/nsChICf1S6kimqDhYDg5+m0AWgB0UJXU
aqjS8dRvyIuIpotE3oQHMsuwVh3+Cu8OJCKMe/vhphIHbp/tf1EXGuvQMwuHFNtNct+6gLjlFXRK
0ehvclRFSF3pHZW5WRtTDOfFzg8sMoYu5rGT0LRjBNfD5QYk/NqlTR5m3vSWaDupiEkNK5gR+G39
hDYhd0Nr5AKwidPjlOHvXtUbrW9X+21eGHE0soNZMcsF4a/vrSmWdd0VBzDDi68lMgvvodigDMPD
Z3mB7p/IbWHCNgfbWD5bfupREaXJXIXw1twJb3mrJqYdlINMkNDMLrGsOIWZkTw9egUYKs6I5wlM
d6y1/hLumMTGpT5nZeEp1pOE5jP6i90KEH3soDspB3OtFhihJVBvtp87CxVj4UxZ7S5Kiv9qNF5T
8JnR6J4orD+PSWjxK0MvZDp+FxU8BY4In8gW1CqYYPgWuuL9byLAtiitfiCgcw06hKJtWtymexTV
ll+JsOmGBKrLewwpjQ7DZmDPIK0bQSJuDIYHmX/fRPgoqC3slwKqXPduUB9GCJdch6osCBIRb4Uc
H97zQLb9vPIFj8ubMUBzPMsu4AFm2GsYExJLHF8wOdH5nMi2cjxGaoU35/lQL2dJpH24YiJKuCS2
+9zQ3X6kYCCMP3uFs2XXtGt5EDzic7Lt2EHHvgTGApWlc/4SMSOngzPM79x3DtLBa/fTDy4OdaSn
LB62uF/d7w3yVFPCZ7Y3Umm1XE31F1wamLiXtmuIxBiTNh21ZpuvIo1m/sL5ezR3YBGIEEfLhoHV
HMfGRYkaFftHDN9NE+T/Kg3+e5cRmIbAkQ/586yuu6JFNPGKzgq4/gtgdpGSp4bK58tx404doT4T
8kxschw84S0Kz/sOgE52nDdyrBzgOt88FNzSEUX41f1M96hLYUgAj/7Myvk4+gns3M2YP0Y4mZgI
fnfXsjjq0tPy9ta8ToQUw9NoSElQxj3hlrDB47ITQYei7vbpmr0JSuSUQhsildbUmqyuQicj6cg4
7NZbjq6Kp7KH6m50LAcowX1U8gvlHRvoC2ZcbW/KFGpdG+2fe0ciDMEp2JxL85dJ9nq2IlnyKBeK
fkmNAtmekA+SYqK6zC4JS15Eh9yaxqmfRxmIRZztI3aJkSOyp5iEXH98dDESWUgKnhrzbSwjreSH
6mO/KD5BqL8/8iuyDMrjpkX+DSK6FjlcgFjlCZUhuYQLnuDY1A0DJlk5WzpHdDAuDnZa0kOdIFh8
fvHuQYcG67V2RtTiaHeCg9dwXKHuR3kARCMMjeEXaOm2JmhaBgquB94YFPKQPwO4efcT003eF9a9
IFDWpSpoaUe8BCjD8WTo7AhdM86+wor+XGyo5hPZvNmw/Zxjs9s4AiencUhijSyvoE4ZA4FIkSy1
3DflDyybJyJXr1bIAZEiXJA5igCtjtMEpBAWQh46b6MfYnI236XhYPScpOmgpVh+sz6y1CMUilUV
5Qzv7ZL+obuznv3C/nTntv93rC4cy12Xi2rKe1qNDio+RGjhLETEOkuul4x6MauXJu0j6U5KKfOv
Zllp30ru0hGWd3QXmTVbXYfdjdxsuvYzgqwHGVre+ogzWHHUj/aKXsQOt/hqmspvvuT9+wnvuW2c
24iEOpSUcD1w+pDl+hj/fItRSZgshvnDO8wqF/gJ6ZVxTyUEDpD5swVoOPkrb67AN8RC/Gun++kX
81T0+5OHnNG870TsuH8bjD8EXWcM6zH8nR2fmbtpJshGizDyxu+FujsOu+s0iQigaL0IlDwB3AA4
ZLa+tfphJiK7FhdYwi3QHj+REWSsP5I4zTKksRFyMQwqM4QGqx1wot0uArUjTKdaLxSAcA/jTgxC
3xStkkB00Mf0qS34hkFhpLQ7e9zfyGCk2xGxY7sc95LQyJJ+/nxnEFLIoaggTQoFyfSP4amjbEM0
QTKBCD9dwGLwZ9q8bgLoPAF6Q9L2GcRDoWk37GcXMTx7LaJuNH+UYYuvUZ7OHSCBNKpOdlXHcwzq
AQvngAzdIuYihq4p9oTbv64lHWWgiF99SY9r32j91DcxrYaePQNAuOQfMTwh39u6owWQVaJQlsLP
AJxQTjQ+QRvzu1U9mVzW10ljso242MZtWX4sgU/ya3RSB0c9vHeiIy3quTIRUu9LpD4y+tR5h13i
HA+mawVumklIOinBm0Ea0rWiHYijoIIela/VFAXsS6q0rVv2vcp8++3wCjeJ25yfNuRtCIagiltt
VlWysfcAryLR9JaYOOfxdv83gRTXxAOGEw1Do88BkIaDfA7DAb3R2b2A96EcPErGgWq8vUM+XAUE
DMVc2cbzsnI66mkhvzYqHhFbwMh8oUiyxM5zr8Z1SPA52dhXADiRIZyEzgnp3VzY5ojoyy45+Go9
fL3f+2VWup9lbnQ+3zG2F7GQ2A/N9Mfcu6apWxLSaFgkr3ThMBntI4qcrxhJ8g0R4TFMDwuy28JA
PWJGE17dGFiV05ueqFnr0sy6iR+BZcVzflf3jfOgfwPo7QTZlZbmsRAlhGFHekG/CGKfQFUWvmJ6
RLQ2LZ5KORberHLsIRiuUrSULFNFC4b7PzLepg3QARCib/2uvIu/asVEtlxf95ZCoPKkBgZwOxp0
4zSjjt2tkHbr0mWKFT5sMs5PwVe5WYqhGUQN5UZsfrQGEaoj4uJrnajlH/bt+2VD7RWU2W30uuXa
57srp6u+fEJJIDRp51Z5DLXtUrF0if7ug15eORRhAgPNBk8TiOB30/KYNvRgRw/irNXPaUm5JClQ
gIR1N6yvYNW7mZxt8IgKQGVVlJ4hPnPfUzDhx2AeAfWKq7a5/twmv7mNY+SEKpS3QISnPNUw6gGC
Bi3I6F4O0UJKnXGrr0Zpf7pgt3o3js0Pqusy5Yn7EFjP5Cd9Nr8Ps3ScO1kCiadU1WZ0kvEdiRBB
tjsIOV0zw217Tg9965FkOkEz9NJB64iAzT8kh38VeO67emcKfpuhnUS2CM1mjQHwDOvje6MQ4pSa
3f5QgrQpAuGoz9uoiQIz3ZI2McMHGQ2sbBcRDNcqwCaHC/IodYAzScjmlITtAo8fEz8yxF8RHXvY
g/3c61K9ZqkbvqB2Ct6gffBBl7PrDyRNyAp5Szu5dIGmRsOt/HlBVsE3WGlfwxOnIvJXzwCBFxFD
zxiv7yZkzKMXe4Urf/VaPQdSQb00xj8iClZbNzW48Zc6e/vWfAnVOcDeTZEPQ2W4P/ynU+umPJkV
QLnAdDUYkp2eR8avB255dbhq/H1XpqZumpI5LtoPfSlCJL5ELhbxBu0WdB8/HwrA6p9VkW5JEPkl
Ul0hYM3UxgKRicenhedZlBFo45nR/UInN0QD/DoCp7Ju41hy7RIv/gZJg/+bRLoPFBS/6OjkSRBM
tSISoTLsA0aFqH7wpibsEFqY5qPA9ktEa+5cl4SEllB7w20TBOdWk6RhzO9keoi6av5i2dHMFY/5
ErzVdCTtJIriCjuaNGOhPUuptLhTBvcTnyEa8odZ5k4v865+ed2oZPOg9GG/0dZxPvYKNc6D16OW
gwNDAo3ESuinuj2g+/TNaAMeUni99DvnFAb1FDitLhqown5jdPBKJAuiEtwBRluWau7xZrvfwlqB
+l2WZteDOd889FID1XFDxKik1etT23y8oc5g/1mwVzkjoxxUb3HSlTgtY+ymjpO7SlR3WbW7nlEl
sVcFZnmTpwZzdvvL7WrFYcwrBtnn7PsUNT+zsbfWaAu410M2aH48lELlow3JQU2S2W1uAKC0pLqz
puoUQgrHuyD78xGcGZCQNjlx6knpPed9Ne3S/5wu5oNkMu/gU6QJbZx090BD+r+/SHVByTtbsm1v
9bf3SewZljq0YnXucW908oQqUJM8s9KDAaBGz8J3Yj36XLZRYvIhHNsWmzzvKRhqeZ//td6yjcyn
i3U52M8lme2+pZhOMdPjVqTOhfIz8zaNy8zCCHfBDtFM8uojJX/oBGSKCZN1SfhsqiCmKq4YjThE
rKh7VSs8FUuIsIHnSTilv0r5P1kNmK4KFtHhjOGHp1zXcc+OcJwWBtH/fHaAp+e0ONRsRBv+4Nd1
AMREB2G62HIHD9Yv6Ds8pG7dJkMe+/OlayChgl09KjpeS3rr4dED9CxrS3TZsyeWm2Ei4fd/uGdO
Ho6MAVA8KopVdLDNG1eQGqONntek6XZDD/VUUMdkEK/BMH+BcsFSAcrnwVjrKpHfjq1ML7SKQcp5
2X+Cz+GLNwKGjUu6aiEVRrgi4Ye7X9MXsqvEmCMo8+UKQe53PT9cZqIY3W0y8LeN42Gze+aHX8DR
Wpt/7cemmwnnoQJtH5j9fm7iY0LopyTumKR08ZQX+ZWAk6XluknMeq1NMeieeguE23WEuNR2Nqm9
BDryqFQmS1ssZmtE+U10sqG2MkRH8ZIsPheYpoLg6zYRQNU30pWeaSsRDlC0yn/hG3TWtY3qxEKj
VDMJGoEmJRqI24jpt0+1cMITnOlDy6Fmmtvqhou8JdcWoepVK6+gcUHP27hjNLbogxq5U8srffq5
jaVAH1Vz99G4NBAdhHk5/yIwiJADa4l98vh1GUC7d8A2cilWK4zgIWLmyoNtb5ofjFfvXOpvqrev
tNHwiXmI+/rnbzI2UH2arwuIwW0g101DTCxDqlqv03dm+l35tdRfvtBSLkEs9Krux2RGtp5Wg5T+
GVS04087LLAbzYpowH/NI1l0hxVt5LM+bs9PKqilZRyzYPEdax5I2UNYiZnA0YB8GrBouHanTda/
pcp9ue0gb3QejhTJKgURi2T69hvZFsEba/FafYwerX2v0ymr9IKAAdD/Gx1MSLo76f9N8w05Wdbc
NNSnUSZYmb8LdpPru5o0VqCKzb6Q8m7XVnwEEgc05rnGNLO27fQpejLgLaUJ8a+tBlHLRkCoAT/L
uJfzGM8aU8K1/sQCa0lXZFaRCETtzaAzCbXLyEtMkbXfNC/BapyZiKY8saciyZcweP2UrdfFu3WN
UsjsDZhgPca0FPwZVVVwB7CIBtJqKjnRrdd8xVkEMwr1n5jfNQ/W3Qe+f2xq7ld87xyaFqPVk2cc
atn4hEr9ewEJRO9MQDn5CWmyKD7M7oGSqjNPZBFefMf4NU2AZwh0q469uHESO9kESVQIMrjKtTgA
ce7cMWrDWXuLBcp8afRFb6SVDI3p0m7ZNJxq6FUqoxLCBd+vgMmH96ry/ogoKijjlxhWIlUaL2ZP
1uri8TH7m1qjzqH7EYTxTtgIQjDwULJqmrOhIymXIwVsHrLXGdRgbc106CjBFBwIIciWVkiIFb3z
mOykKBPlfE89PErUQsT+XmMuNkI2OXkjk5Ox+3g0ojhRFKYBO8RpP4xptDAHDONjrxTW4I6YWTnK
zU+q8r3pnUT1xNR1QBMhi6t+WY+noQtxTmBr9Tm/ef5Z9l7/lKfIXM0mtsWr27CLJNbQpF8U88zV
MZpRXsqlW+JC8s+V0DsQ2NuaeeMY0VFNSp3NtB6X4pqjbjc8DcgFlNGpltmrSm1K18MYtPd5DW5M
M8EFtUFslMAa4TMH1b3DPH0xds5z5QVZxVdG9Q+NZZGnaQZ63NKf3n26OjrhB7rB0ytcAr8JCEwY
TmrcWT8A+biPornTnx4UO8eqCk66qUUUDAJabR119ueRKXzBdLa5v2GvW3v+yRpG3uFUt/AUrJRy
Ixv+L71KLV5lYcXq3dtVZwfeyyXUlS7r8u39Y6fHGo9cXh5hjgpdBeGUL35I3+Nwq3vlxn5yoTkE
ih1lKvbB6tzOu5jaPmBcdq7qm7GDfXxHxZRCfWIASeDOTBXS8I3UtAwC0VXJ5ytxvfDE5FaIbjbm
tL79tEOA3nzQ3XLfkh7EPUv+lPl6iv8r4EYoNxcb30y5Z9thRn2tp6NupRRtaBXKtIhBY1wzs2Dp
kQ1pGL27sXnkSfj+IWGscS+3YDFBEy33d9Ry6E5uc5BMOSnyIF3DRjgdVzZCKwkXV1fWMt+pFOeW
PW2qKrvzIYO++oA2sJhkhNkQ598yFmLvTMDx6cBZTQ6lYqnNUfziLTODGgiUGD5rmAGhewGovpJv
1IJXHveoaotQx3KbAXC2Q7cZUMGdpcJiz2tnW6repFWcAdgc07ESMpqymhO3+Ti7NfcCNZ1gi0R/
EanYfYG/yZ77Wq2jIkpYOEkG1uiUw3Xk99nmg9np5iqHarYj3XsyFzuLssActNMbQ5WRNEj645M4
qgpFYj4uAG95rHhqdH0mX0ogogUXxh9hizNJIwNlZuScscg2wt5rcgjWjljnlNraUKzpNjnQnJAw
jJxrGrvsbdJpHA4QPYnnLukmoBFcnPe4fq4c37WlRebn2Xmw/W7B0qX/L63ffkUjHJ0YivHSPk9r
hKuowfEy1OstAJPVlbfHOSkK9z5HDjHjhefZ1Bia+r7RjOHqZ0bKpBZReMWoK4QvB4pDWO7w6TYV
pEbJLjkLnPU6uI0eojfT3XVN+XkRXdRKGXsix46/W5cqK8Mbwo2+3llnXRf48LnfIiAtn+UBcmwA
TGNs0I/gjDMrfhEQw6iq4kjQbkXGSxyskHziYiRKEx9G3vX0YbB8b4qx33JNCZoEcQK73MeewST1
SdJNNEXS0c4WC9N+HUNZZpEOySgUEMVOKnnDL2hB0GymiyUeVfT6lUJaQsKAK6OJld6XWOHvUPev
/ZeY1gyxLWfeD66+1ZXBBEKgeM2JrE26UoabBn3KGgHrc8B0F6V+TcgTthyZYpHuG/9dHolwijUv
3hJekM5tryZgwVBcInEAVd6NjcyypR1o8km16IUam6Afps7tedLY5H6xueSk275547Juf94HcrLv
J9P1rTV3VqiPnOhncu12lKFE5seRv4YOo0CAEYMjktDzi8dZQ32t67fs5asZqNAXjNM6T3j8pO/U
v/2g1VFARuC0+lOq8ozJrh7PyAjnF0+6ySVic8p452g4WCKIs9/wjy1Y4PRq5EfqRj+aHyx6lvLt
tyH0hu50RhuW+v9yChrT+qsAkXbNXPfM2EGjs0Bd8xGiGHlsWzL7F7Jk/ROxqgxSgtfBZtJtVQES
N8PMqPEAYxL3rLdTwhnaQFVUXmTjNG7wIM/Te5yl1lQikbYWmoXoZupNKvjCzVWQu4+Vj1zxRxIX
dSI7WqJleZWsddwxVwIwe0NGtM4TmmRDMHqI41DR9RvxHsjS0DkAIKYnMl2P3qM1NSRh84HydRJ7
keu1Yr7ILp1G9dJBiaArA6Zrgu9oF/K8HFPjtV9FK+bKnmGnEccP1UuzecienZs9fIui1V8KadIs
EmBXNEkawS8cmlY9ny98QoTdrpIBLOrMA86PU27QOIfFb+pEr8+vUfgZu3fhXa0Tc7A1lHZU+ZLc
xxTb2T8thzgOjBQFQM9bsiyURCVyh4iCRrK0BVmdMuKdYJRZdQcRYuFF3TfiPccprgmqpEtJE4AF
pcXNtw1AZnfwqyaAoXKi0siCCg7rb6SsDffgreoDb1DftM59AqKOGJVtsf365z9Px0UbMOYZdt4N
ImPnCmfrolvuqXElMHAH7s6DSSLTh0LYV7/VF65x3e4j+/+qFH60U4sVRR9bOajUdSRabolnPVxU
+5/0cLKdyGwapADA1ub8RclWNnb7hAUJBSQwnH0IADEkSotosibeV05BDl36wiUNS4Pt5vahefpM
bCz3N25YUKeixKHQFJn00JNA0hgL6lPW5q0DDHsG+RbRK8Lst/Ofmest0x1zuI8PmZ606clVnUIn
hkiO8WNr4n3TpxC0n6h4mXA+cEN+NXgWsaZ9YCoi4MGCj9pcANEwvp8wUK0pYfhLgmW4VLiiDdG2
7un/M3PAVdlTmkefiUQaADqrafJBDqTHgdHV/ZFkKXQ+Eb8+/8xtfUDUdwMQd/fSr0bwH6wXb7gG
Zpvx8mozE1kGiQxi0+zaL5uPSAebLeDpX2FarUSIyBN+Ytm8I/dn8KY+R5dVp45eVZEftOTLvoOf
I3P4ukfXDW1Zu7t3yrUZfaC9lS2Kzc7MXq304FNkVBfbs0G8X2mvvGFkq5VnuThoqUYc4Z9OOo3H
86p+ULNxZ0P2UKTszdHRDKSXtmjkpul9nOtROlGVz8vDOKkFeuwipOFmPA3jFeCRna7PGezLr0Rd
KRNdRlsz5AktVaWOvOsYe8c88TEwSvtSXm4Jzlj3Q9jceLq9OFG414/EGHxCc+0ulhx9rGB0XN/z
EVA07xgO+1tSbYoXQ1REk6wO+XbqW9Yk+KP3rBvs3H4e7E9xJV9qRtlcmU8/l6ygbYGHTQx24kI0
BoPp/elJN4AjrqmJJKLXCe1n++ISQVClkEa7Tu9rjo3xYyrKk1XnpRnPdy6eTNHzt8wmp2QvViUo
jiYEHBcwyjDmFNGIxxduWYjqbqTTYuX/AzrYKz/+crostlqVHN3O6QIKBQJB7Uj1qzO8/7slsCUd
g1AvvTG06Br6VRlnEAQ+2usPdPZw9+94exa6pGaGDj/e5PaK7L0mi54YEIfuk4yfph+41CaOp+aJ
UGphU2Mh2YteJeXKjC0f5eXM2SjRqDMeEyOlAlA9c02oFn9NnSjGEMOmujm9cyNAxrhs/Vk0nE6x
D8x6b4rtoi9n0SmuGFdMh4n0EQJDsRyELcdz9P2+W6Sfbsr/db8QsmawB5vX7NbmaNrATg7Fibbt
TJvISRq3WV61upcCX+Il/tGl3H7AzSwSfsXziQGZr9ULm8KffbdgcialH1YYLgAA8KVzHKrReZOu
ia+qAOYs62dtNgAuULcJnVFIur6LFl5bqZFgxZDbImQpaq/Y5zXW7DKG7s+bmD+UB2xPcPeufbEe
cjuLDx9WsOPneiG3WGP+F8SKT+3ZNt0upJGrwZhfZamNJz5cqMkl/rSooGJbHA5iE4+w5dxC9IXL
xa8b5fJ0M7w9yYpKz6jAPYhL0GWxNP3k8DckS8UewyELogPu4zzg3CRhwa27YJ+NLcfNggFb0Say
vNdWCJ/HAxxV8SAkjzu4cSEa9j6XdVSP9ndJ2dAuvmgQ1Esn3RS3Qd432uGU8kCRlql4m+3zkN5i
/fUKwt8alvGiWolPLKm5zUj8R2JCowzH0JUy7wK6JwJoWXasRD2Qx3aRIHnbj7l45TrnB7Fs8DKb
z4TMbxdVTx5Z168Y2eAyYIIk85raPOe4PYGK10e+UlU2X6KFT2ybUN99P+zXToxIHEr9usyaI2cK
X6n5867IftEb+FpqFmkCraRvNX+F4+qEysQi+NKCjo1bK+GUFr3T8KOV5zfKYjyedGtlr8dSB5Ua
XzlUOHf1Mf8b5pvdlY6gB5vVVl2RZyZaqXzdmtgQ5dvu7vIoh12yGeUIILIYs8IdcKQUi+I/VVy5
vq2WlYCmnccEjWeNh50PcApyUYtPwlQofOdcPVE8vI6/yvzajqVLLKd4y+au1WuEJoAw889Fyeng
I3I2woJJTxjRycksEV1WtlC8LoeCG7aMBKE35W1OgvxfZkVjAB3BuZjPDRglyxWC5hVz8OASRE/U
/zP7pBtEM0PNAhh5jJJE2cN5GE+k6U511yDy4eZfHI6p3fo5DaqQQU93Yjqd9Tozv7zQV2PiRV92
QV2QnpylWdsXBFJnuI8RH64cSWDukvSRP3I675sJIHEtXb8X/04H8FjCpkZEZGKPiw+TephbQl5i
jXOioZ3IrWp1ih4NCpcSE1EKjz6xGBsFzwmlOYHSOwXwruemW9hozz7dmwNUK2Elh/MMvCw0aeTx
R5XlWdiPsBJKNoZGhgkSMXQojDkp2nIdC2mKMTiRdcgGu9NQ3ztuaLwYUvUyOiQJPTW/HXYJY69p
sKaC412bQyVwS3EEhKDYtPkm7w6O4x+lVJTYeIe6uqco5YTV7St664DkZMmriXxvLYp4uMap9CMo
jG/YLMVTbnGUMklKTo9qCLVLJx91JLR6qm4XaRInm6qbHutEIWZIFP0FAgBH79Gth6LBM0gTh7+M
wmrI6V4aR1R5d2DlFvzZP2eYLAJxCVrkrfViXe4gFWeYv0XD9N99xGlO1HcCIqPgFNrugQJHJrnF
QNp4nQgxptoMY02IE75DpeM2J93wOUXUkDD3NyMypAD+vAakn2PacdJv/RfOf6ckhuwMhXTwkL8e
caNMuwKdPHQqKf+PAim3y8QJidb3/nCJikSU0uM0rl8iyqSHRLoUCRe/Pc3iWSw2N36VC2tjnNI9
EDxHgJwTUbKuf8m9F51uFC/cNjhP1aMcQ/nU5I5SwvknjXsFfSjA1p76WkcTNugtDqsf48qjtTRo
TlzPTXzV2Yyd0vTQMMdJTUfa1d4gZuoQQTfQWQX/uxnkXjbtjtrhr4R/Ovj7VePJEIBmhZewEZrF
AmXbdwcwEQ1pCCn1GIA1HhViazuYZIRuKLjfwOPU0avpkC7mVQWEvUPCDXBywuwPfvZJMkhef8QL
3KTCn4HJ4hSE1fCvbYXNyyWRDWeXTCOGf8Vzpkeq18b4Ogpzk1vIeWaXmkT2pXP3MpeJpN9c3Hzu
D7uCV15A5g4zdlYTvlVHk6qKGf76gXZlYAdZ39mikayNhcMfv6r0rVF9qydP7xH++5ndAD10Tswi
NWTXwdZvpBLs1NxWSYCwVrQeWxuYOzuzfgkwRyBmqB4NCSdTiOnAzyZd9BoldIDtdd4xtEiV0wEt
bUfTkVSXnYRXgI067rswhKbrKUJNLxKL2EnDJxxF+E8FmByl41nyW12E/C/TKSeO7Nc9U4LefBWo
CJmKSvJvb7k5+4uU5IgFZKRRurt0u1bHGic9ieREA/5fNAI3yB1fXZzbl1uLRVhAA8ckY+lGOXlf
M+hwJl6CkWG9wPS4p7BEgaBYSAD5kHgHnudXZiocbcNwUbFauf7+YKy941/Ige2d19KmwmX3EWoS
zHSOBYtOEyMaXwabyyE5UNMS8H6I3btpxkyFkajDFgalEgIKUYE06RDeRTYZ23bPedYYidssUTlh
/PXjywE4/Uc7TXo4pgjqJ5OLTosPhuFQqUqE4SwxO0BxZhON1J/rM/MY60tb4Cjt5RDdDO4CcSQl
TkT7pocJdSylcbpLBuMzW0lc7rq4AtlafJnFcuuf1yCP765UapPZkYZLsNyjDJ4/ChKXyrwO4X8s
zh/jV2Ki/Nsi6A+u2G9MLRTjD8mYgubT+J90XqbxN2wBvWx6PclDpm3nxKD9qQMa0aN1wkKH7Q57
TM6GyKLbOYuVbop/bP6giiwKGJHtnGvkCU16Nk46xygQX+sDU2FnkBQCDVBXelj3hF9oa82wH5nZ
XrtVnT+kv3FC9iA1cjcK6h2Bjj/sZNoJ5OTCOYUyq46IosXUHBrCAS/cTtwRJH0kuEQ2inC8/q2l
cP9FkzrJjtWF7mD3K8SQorxjA15iSRyF/eHvSlXQeEmwZ6vvkUzGECu1XAkeqEVStjC4rAhvQU1N
uWu9jEqWPhlxYM3TWjBqsRTkK7qaSAzUr6pEERPrYcYfPbq75T+2meCih42vk1W3qz8yza90xVMn
E68WcySCVwRkPjqwOfsc4Jg5yApVZ/DD3s8brn/z/3reIDmiSDh1bKHGI6RtF8Zo/KDmtZGH9IU/
FasQlb82G5vKtoUM0T1osOscJw1IJ/12lCLFbdU1GwcZoSkl4BLK2SKs590m9X9sG0N8QNY5eUAL
iumqdAr1uo0Zin44j8yQ/aXuSa64Kz69e86E1rLBPimh3mLK+0IgBovl3/skg7TqGPK8AY2j0dgt
Q7MZmVIU0Gun8OSf6eNC7/Nk3h9U1QxvbFLqg61Jiy0yEmwGvkPQxVY8dW/7rPPBqorQetIRywcm
xIdzu3mLJ0EuMsuTP/GN33KyknfdLNTHxwScNC9WrgC6S4h8s+nnNcYQ0ga96JE/+EvXK2pfT92L
6PMnj6F+7B9lgZn4lqSkcTFXWU3krsqGXStxtbKsMNtuNPs7RABq8B/cX9yXL6RwRFyIOpm7va+q
asVEmKhtovA9qnobe9O6KQdgR1qHSk+yf4dSAfbxBTRFL197yfjiMF7v9c247+jRyVla2cvb6YTA
JCK5woHMbAauYxgdZfDivWZxvE7Rqv1tTFQCmz6KyErsUtX86iP6OQKtGn900CjXUcG5MthXvT3f
LVf5Le5l4oBucmhRLXopzPDlViT6C3TyjzkCpEVTJ2n2aMKyDq4hD9yvKNm6OnFsowf1NFkcHaMo
wzACIRk6FBCNf21WoRC95RuZZKLqQ0vOxV1ZJovx+j6Jy4cWqlwmOmJyxzoPoeLevKVc6NbimzNO
8LIjhIH06K0xwzptreMA6APZaB+1QcelMOTXDNHjfbCJqFnQhI69UIOEcKgNTn2vMLw8LiaZyR5q
bZk+fT6bADpn++e4Y1b0QJVk2xZPXxziM7IBDYXOSBJViO/FdGl32D4CrDBfzqixIGhZbytGKb1w
fhyX7Qot5UOyfBTfR8iIGmAkProFzHPzrfXOjKtOwHxDfquWg4zjwgFLErjgPfp3wgakOpLDmjQg
SKEQ6quIsWP2tRho0gBBwq6uAJHJ4RqADEKwMnKL1vDueUz3C1R000Ugy2FK5XN3WOsqDZpcuTW6
tTN7551/N2JA4fso5wxg/wuf6VtA5Pbi+ISrj3dTgJLJ4tPQpRwqFmwcjhogP6UtXwRFjvMzMyIk
luEMY8EqiA8xQvsNooutBmGnI2K7pvLTLlgZCHgQKp2nHa1KGUbtvdKLDcoI/QdgWUpCYnN2mTUA
aNksCLWJJhhsFelVHS4BYEO4GNy53/UJa0KYmCbo5T1DDRQ8jMGoGPEWpKPAeNovsMqAwwCPeDW4
DvM0iF9yupjCU7+iFdnZgLxK14x+uNX3VWXcMgzus5QfSMVb96wLJZbzHmyRIKV6MlZCsqS3swc1
wtzKGbm97WqG3eRDv3c449qplyvxqjb4G6xLBu2hQe1I0RZIX2ZZ2mUOc7LB28IyHbY3X2UXYZPA
i7fa6Xm+bOaE+agrorLYLWmEhX22/u98WPpmZ0y8v4uoJs4svxPn4M7Bpe6C6ONJ2sZpJJALmnAQ
Pl9XNrv2V9KUYCJUu0ouGEPAZLxbI0VnafkVMAxGK7T/M24aihsIQgH4UlugHwX8dqiXloeIkb9h
lCoHeTgZ+0njccpNdkO+YmOUdCaItVTfaVdWQZzYpydlF1Loyzo/EwZZ+fAzJkIgUN+DQfYQCa7j
ijzlHDlVN/tJ9RJY3JiUNzZzzyxO3RZKASK0ybq3K32M84KpFFVShmnZ8vxwUE9/6nnWkYghwS5a
3r/ooMguRdYoi2jaJmED/aklD6KsWYOE4S7F3+C0rRkBtAdnWCLVhIFVRxobuaT2he96AaKFjhl+
p6QKfW1CiJr+cuI8bnuUBm6AXSrkOK0sLmKrZA2MMMRGMXwKRpC6AqjspmFXJApbvJRF0ifjvIN0
STsTmDEsjNoTVuNAYzLLaXHc4E1rTRIJh81gPVoFYQbze4kj42yyC4CJ8DdRsAwO+2XFyPbpvvfn
EBe0ebxzK7Hi5ErLbke3ezhGi3p2D4gaWhxjWmuKWlURzF0cO6kTfWRoGQvayJTlCfeuWNF/wspb
ZME7Hurkrlwg95fFr3GhPuwSNWP5Q6D6f4i2xpeVoqsVmPyOlvPLVWzMmdvsvXMQDxm8bF12jX1s
s7OauA+UafAtENloo0F54NVaOwHFGvW0PNR70v0x/gMPdIUllSrWrlMJ3g/9cWksL0WQ7YmcXdfh
Ku9dqqON+Z26sIvxq7s5noPC9JkA9wvN/0QwjdQAhb1Nak2ODVx6vBwJx8ieZyrpWWE7Mp+LvNTH
IWhNqS7urrDfBUjQXr28WVNJxdbuc1dn7O7mzdkNovHFpkiKQqIXXu/5wGosm/6vFQNG8QPj1z0T
cjYLgMyC3VyYGjNWCqWzbDNEZs6B+Wq8iCLwbp1FUwNp00Sw2PYXrM0JV+wgepokT4XWUFWN0nHr
AODu36hRTOZCbgdXCRWHgPR7ghsbE/CtJbVcvshR3+ed8N/p5znf5LHXnlyFBnNYmjVFw6IotV76
usQv0c5HwyUZXqOSIpnw60YXjv1opHmdN0mP7zXHaUouLy9v0d2ZqT8c7IXMEpkGiNJnsPF05FIR
tEFey7lgUQai5chqeWs0xyTe4ZYqUoWdwoqpFCp4rvzmfNpNo267ECSfBMX1ato1sfzaKU3obpxD
qS5yOwg8Wr/eOdnZk7Gv74dfshWdUE6CKVuHTQm+Iwql3evo4DkCg5GPQKQ50GTDJ0O8aIKVXPMI
QIkAbV0+FzlFRTv+Vw5HTSlCNr/sb3jo8FmI8RfyBaPqtyvK8q/7bxQni0+t7mfjV2tGLYO0GMA3
0vgIaKsGvWFr72tk3C5tE9gCGZd5eDWQ4275V5djGCBFX+eRTNC42Liqg1OayA7LJJo82+zfsI1n
j7aicjbevJDQFYxz2QsBHlWjbmRYBY75Rb7CVZVl4QUffZvr80BM255JSEk1QzKt2Y46deHKAxSS
7ZHyF6tx4B0V3Mw9vFxEx8brHz6X01x+Qo+uh6JyNPiKDZYOF8F0I5bbgxyxoBlLFRbJnnE3S/zy
vvPTNjs+/+TXxs2QFB1qjArY4m8s8ZDMAqDt3DFu4ZyUij81tHSx177rDGdPffMgDHdrgDTmT0Pe
uVwUXmf0MPiJq9bL10c0Y1GQr8jGR86SSECaT+wEDo19TvxvVYs3FaSLymCL9GEpMyDrtPwdKSDv
vYDDNOu0hJhRqZgKU6eF72bePC6u7OZg4/3alI5XQSRFRMABFsYuJD9rxlByUoYforns1mjf30ny
V99zeCWlOToSI8UBJF2UK75pk3un6mRpwTe9NLVNyqcIzDW2nNZKlxpnTx+qqQPLOYbxg2AwROui
HcbiDnzS54MvsBCBrvOU3PPlKXv+1/+6WDRhL7I0b2dDEZoGtCiTZSLc/frPVumFoLcNlQzu/7Ru
Ze8ZarEoXSD8T5lSCCedcWOVOPA/gL2tudrxBmGga6apyXFm6uNpurVA6ATamgHWyaWRLH6e+fRG
/eoQOQZus5bxJJFu5V5Hxtb+uf/qjNEsZ7UTPcmtpWd6SVrulVBtLucdugGKOeSdUSPLuhpEWcZt
5diUwVgFIb70v4bSJLvlfqHjFPrcGWCkclZ11atgE02sCn6bIyGVJZngWyEhH/wej8tQYJDrDL1Y
rdolH8jxaqL77oAf4EfTC3FD5RvUYDQ5KrgJqgFqHp1fgx9BPjYm8B/LHmDvITbTssjHxVQtxBG3
g55SxbvAqu1kezZ6bPiYy8XsvjntkE2KxQe8F4uHehBWohyTl81/sU0XrbVA9rS/1g7Kxz5gYTOY
cXhHntu8KlahNsJpSF/qDAQUMHXfKreXlrYC/MaGlDomHdx/JRf5O0ZLLcvzFnvZvVCESE/9VHJR
uBq8xKrVPSJsoR3J1uB19SOHnA6H9VukQFg0prYQnsJ1H/iQdBVT1NOg3+nqJVOwHUQ3TW2EeWqt
3TiVeZoblg0oC+9MhHfoI8t3vfTFdvetARmR5njBbEgUCFsK9ZGcnAfSzQsuF6MZjOOtgcecgsxN
nXx9VbncfdWjmH3flctjrn9TNxp/KmIj2DGBanMjZCIYPI8iD0Ra616r/hnA6IZTm5Lb9pAM/Vpw
1OrLBMvEZ3EauxTsC5bPUzroIxRaFHqw8ODBe95HrL9jTIi91zjqAxaoeHHw82u0URqP+apa7DJU
YUpjyl8svqV25rDn9A/yLVpfIQ/UCSnsx2b1ru6o4Wf0aXqjA4rM0ga6r9Lnvu9PKQOasnDeQbMD
CriA1goQ1aAKV/mDjuA8c3h9L1HvaD2KQF8VRwbtDP9YIuueHmtE4ac/bQUHnLWSJeO6RN8YtnDE
LMCmP8EYtN48avcGtjhDwYtN867aZiBcphlfA3UPsXR6RZl81Dn2tvFKd659LQX2sLdZe9qZEHTp
0awZhicFnHGeaeksFlnQswhjugUAzFcl68Mwa932TQ/TN5hmD4rOi3YRrstfPu+fPHmrBCeCH6wM
naAS+CelbeEx9eN7JqoiNM1KmKNFy/NW3bYYbuHPXBg/T08ZahhR2DYVA+yODZjAL9LQ0hlH0fMA
SzH1kX6yHVl9LX0MfGb4I/Uadeq9xP6EBHJ5A74+FE2PbCuN7UiQKk7LCiW/sveHBgiCB4rPQ+Tu
uIrPXOHNXcvtVpSy5S3+gWb9Gi/6lgTMfSC6YdZdZLpLGZMN4q8y2KDaKKGNIu4NpH7uJLeg96pE
WDaVbOqbtuQwkw6tRIMWh/U5lA3RD9WIaYuC/KRCwTRT93tMCvORCOqMhjGE1OtK9o3+2SnrS7oe
djpcyQxKlH+WkCjB+3Dag2g22PgEUQHUPeZJ1Z7hcgOZ0wg+XwXBqDfa2FRqRDGb+/c1gCUiG9ac
DC7SuEMTy8CB9D59MiIQM6wNaykHsC0ztE1JHOlwJV2l0AxXTFAi7D4kkMuPWRIxUlJDTQBThBw3
YEmb1kJmIA0wZw+KNxwxcY6NeET8UtmU/NgCM08VNiAZ5cYh+7gbo2LaKrjUiY0icWgV3dCofjTb
H79I0tiA9m6hMvPOlwUDzNS+c6CK44KX1MeL4CBfMot58pUxw37mYk5HMaOzfbh8jEeoFYUDecUa
zeuPxGfvoMVb9NV80BKU9lc1Bt/Dl3XkUYMwceG/yC5xP5vzWVKUj5tE4NjhIR6WvLCBFQAVLCf+
LbDKNKvXAVpiC280JVf/0xO8ZksGpXleoMbRnaP8Nrq8LfS3NFh3F18ZJtn+Ko2XyDdFC5q/E4g1
8GTw1J/GJgc3rcZwRZPgFseyTCOVNZfVS70mV8zKBDcc0yAbP1Y3b/OS63ZCK0lULaBhueuAZIP9
kLTlALxK2R+qNvz50CX/4M/TKH3zCrZZ23sK4a4oj3UoeFuOFT5HDCZtV2X9+RhS9Wto0RNgU9tu
dAYjQkIJnXA1dNIt2rY4QDjWiruV54n4/kghzWsnMi1DB8ermajxZ3/X2m7xYX5urUoNOa+Vn5Uc
tVeGxOuLRewakMDYFhomxuz52+98BG3ntMipjG1XnabqMAp0SZhcKd+BogMu7CIQC4DdVuWimaW5
IPormXPiYg+FLARBNKAJMFUKkVDd6W64FPHHybCh6TjbTIohD6DujZIfo3qOdIU7BMLv1pyFpLoK
NyKbQ+qluI4VQ1MvfY+udH/lgWUTjsuA74VytwgtrcZisot7BlXg3HgHyrisKKQiAHBzgSb1nu/U
kEjMM/TJ+D/vT6qwJ2imTdOr8QLrCoakATLoxatTCrCkSyL02UbgwreneKpG05sA7o5SdlhsVQmU
DMMm/xhBuZV6prsAj35nS5ra6l8A3mduDCuIEsikJ+H+s5hNvhj985BZnWH/i2Xf8Aq/CTPlG5SI
U8ISwo/YbRUxiI4hGUKHTIpgGET+ckZub+W/DDt+2LYEdsF/gIAdHhFr46qvwgyTe6MoSF+NG2gO
13JghoC8ao1iFwD80BxKIE5faALmvPOtKwHW22mp+R3LriaZ4zB9QyM0p+VbCGBjVj0CbTpz+dRF
olJC6CX2habYOrryneGYhlWPZstuz437lshWQXmDJp2zEc5t+V0lHG2CMEDdZv91XQqVN4MGsR3D
YBTEumwaI9nhaLnxyAyzNkUgszxMw5c5zvFddJmwcSZj9B+RCYdG3z26f4ZSbsNE57lLDM7pg9fu
s1//+9Ce17ZCC7p33VLRIssdJnt98+5iVws88pi7nmoAFJcr+YTU+OZXPmxLTFi4W3t7bSfhiEbG
yzm0IfC3JWZbUcOSwBZhC6VzzN9kGOOMtS5+avHgpE7/BRf+UwRaYezNrZ4sIt6m5m79QSyuXarH
lG4ezBZwooqyBYST5KD2Y/psrVEf5IaEBY1c31YSpxEWCKrXH8Nw7Irk0dwaK2e5Bd3gl6j5Ll5N
xtkMipMfek1jGJ/WvZQQT69RvZEJb2L5bBBZZtWz6H9iD33eT7tVNdimhQpOYPN8puoM/rQU1d6g
TSrYthhQbWOsvp8o5UDiB3c1AFLSp6+0l6I35EArIDOT4DljXTrTbWyT98jKr0lHl/qvLGEGP6pQ
dQ/lBtt+WSiO/HxzgZzV5n7bDW/uhfxIhCZpsjnDZ0ux8mgu5iQK8vZwyGyaI+a5x9nOdANh+brY
t6zGAjAMMh3LfS4iZy2yt+aHhJdNEORItdHa+WzhZMbwRRNSA/a53RU9A1cHY+igd6k5JDnZsAk4
GKR1UMjTwD4QM7aI5gCFZXO1HTO4hHhdP7wGvBTLz6HsFlYwS+a5PDFLszgu0arc1htmOqaRLeAc
9Ud7XnINttqH93x0ta4ryFk7Gt25Q/a+vWiSShT8//KAuvdgTFNsIgeMwdFfG7rauKQkq8AKLc8b
6C7FLv9RL52AUYR14mJIStacVOXxeqy05KFl7AFYemFYuQHNdQTAxehJqz3kYlyiLecSaLTmpz91
NiOxw5DFY/eqY2j9+ssA2JLI9a46avHTf6lqZFyMfJS5La3+UeJFucCWivXHcQz4V5pzKJ0+VvNw
+Pj0dqFfEq71wG5GrYEtnVjyhkKn0suL0jhUW8k02F5nPGOU9Zond5UFYt2Bh34fMAmnDZrmrXCU
n9BuYNNRyvCpAgbOUVZLlEnDf198XourlISkrrLTU8OSTKpkfs2e+6XhkY/LMCO9rwkj0EfRUZuQ
S95gf1ZmAoviQH1snqc9dcbBw9cPDFgi6jetQTJaDAvEbR5H3XwfDYDb0pXr9WHPC7RH92wY81MP
LqbmqbIB5eEJpFiwhz8cQZQCXX7PRPwv+Jte3vSQ5q0fXebQTQgHpr31TrOXK0g2fM9sCuJ8DUPa
nwvFimQLFAV2fxTVQbUC2QRIOLf6sdmZVZvWhXMz5U/u4CYSkiOmHl7hWp8KCsakzA2Xv7aQ6hp2
j76ySeqICh2cW5HHSwiEP5VuBJWQI8jp1+sPHagZ9zPQeMeZkVntuJQMgucIWeYqysOiV0wEkUOU
SA2UA6LDKBdefNLAjeFPL+pPh6nnYyhYqMaydMt3nL5AYgqlhUXanq48/qZN3UTpNbVBy0qNdoXz
PdaFDMIwRw9+5fbb441C5AW15MI4Uc8vHWWIL3PS+gg50ZgDd5671Ixn1rBlU8Z6kSUAJpawzys0
SWE34X+bDNeCxOwPkGytcDohdN17mjPqKE9a4UovtaBMI0eXC/edpyRLfT4mhjo7LX2n8NFIyxDn
U2NLLIDX+F5bDbdO06Zx1AsTh70mtxUXMAhpnJk4gN6Dtzjo3nL7rtDglHWxYt+cYWEm9yH1dtnZ
w4ubT2zir+4yyMcsxlrWjbQ6UCZyG3WIUbuaRfOGWt0OQCVFGoypC5TxfgsMJlDZm+ZgDk04ZWNP
drx3T5eBBSMapL3wj4QzDmSI9cH0QyTg0EX5pRfmJC5mXxmIaM/gOBCosR2qu44SsXCEhS/tLxaK
ukBYSTD9IGvP4jjw9vjy68I4BXHajdB1gqOt3xqgFlf3uTkwhrjaHmLu7PV/zVIfogLV/QjKUCZQ
EJhuWBU2iMznfU6honcbgtkYHe/0K3rkczkmijh8mlBA7AmQN2VMDIy1aRRu8FqFoK7HIr/pVmMy
C24m6E8WY+kZZSheQi+0zlrc3eMhjnC0pGnTVORnZe4HJCSUDTZIUNJchq6/pdL/8ib3DkdtxU1R
KjiDMAQhA8pO46YGcG5Rjm0ASHMwX0lN3ZMp5rRcvZMUdXHjXU+b7/pKyll7WSS3qnbpeo79aRm/
RJyvPGeHLzkPGgOgArcrE71eHJJEVn/EP1AuUbcRe64wK+U/xFLxsz0ag4wpxqd84m52DqpwMsBg
oMs98xI9WbSa1SBBKSBpKnhhYvJRmjF0JTRlxWEXXr2B++ilmX+I3DCipw06dVMKT02idGkhIbdS
WXQE2xBTGat0+9zly02AkOlDJZ/JvnSVLISrO/6jU4gyPpFbz3z0zo2u9k25lqJTIBC+oyE9Hh1k
eF3CHvlYVyoyA0BO2IqkAgtnW9Y5wme/gQdG0RlfXohVf7DE2ImS/L2UEKg55feB2SGfIc+AEP0t
XcLoh7j9DQJ9pJBUS/N+14VBQwnqIDvfyDVCdtjUUgDgLkXpnbpMX5ObNiPm5kiPXUFDA9vFBZ8K
pleVfxv2/m51xfwhymmvkbG89kLCwxLNj9b4FPapPs97k5AV2TBqyyQzNA3SnAGqJTwliy4f6tdB
yhIQfDXLM7zE6sK0OEswYRsdBQRqW1Oo5zlHXZJa9l8fhZZsu4I1gvYZrZnMO5lbFzeEiG0rOIq8
8mkqHBIRPZaiPFsBXIveo/HX0gbkUL2ueVVGc76Hplx8Yao7UV7qP0oVsUYiM0qZN+wS0mz96seW
4q1Mkqs+eZD2Wakjg55Q6XyuBJMhEGdqqFPQhoxoR/HcB4nXDhZrYBOYy7u7G1M6Bmqm/cEpmSsK
a8S2JjecXFuZ02F1Temdc52Y0cp8A7MwscJtOtKe714aaGZjeUn8P6pS1QykkWyuS8vuUNTWus2X
/87cQZigcDJhMb7pPvB0TcovRcmz7plSfSVyIgbYdH5z2Rk4nQjkXLtD49Ow0C2pAtA+kpTk/gZi
/1hWTJQCJTGRzHQEB1Zq1PsSk0cnasB/53nrcNVSRMmfh6l/yST12ZABPso7qFQ/jr55w7Fbdpxt
ErRyf1a9Q9VbJMBSsXi5rIai+N/vcBbrHTN8VP84oFqw/qC28TFh4yGcTAALf/pEFS4ssEUqoEht
vsBfCCU+zoDcEBDxQ2cAEEy4yL5RjvhSvguERz1jWresqO5Mp6LtQPQQ4/cJ73SjKJnmfEgKRfhJ
9mM9tYV5Ho9EfnQuupqfJMtQPNlQYnQFIvPnxrAAC8GogHnL54pCnB2jbLs7qA1TXSDM0FxGooR0
M97ZhteLeAZMFbN5WOzoj8CsI5LcUib+RwGzMsN0mUqIFI++a2fpaf250+xvd18zNQMf1DnFX7SL
j6FKuY5spZqI2qq7tA4YFxk11l7ek3iCkzFdWea0spn87DQCSfLgsal4gn4UctZz1PJX5E6NIvqg
HWj2dPmEhbHTAuNwCpRbExFHgpvt7q5rQcxeq3KPnljHlBAAZaV/9ILKu0acb4eaW70C0wI4Lpjf
ECv/bV+asQHdqNBYneVPs7qyyPNjSMR1x9LM0vw/8ksZceLBKDZtzGrGpY4HlgoPJsrA2EuknPEs
PeWDGGBxS+PpEwlCVxe4l1DkDPfBg/L8tanbKqemmDRflkqnSZWHyEWmF4hTe53tFVdYNHbf/jOQ
c/lcWtT5tVWK30HstupFzREBCXDzZM/FBpFrH5gEo/m31omtZxoiQQjFffTYZrfwLgNzeMMd52Zb
PkoRDMenJdZdRL9igjdy2VU560ppGvW/w47uYIW+BUOTgDb99F80XGJ795lgD6QEa6k9MXARI13G
uRnI3/tM2C/qwgA5LkvqMpgzCHFcNvObdNasCVOjwR67sRWwWNsLXEo1ZxJ+/G191GS1P8SVk15/
ibOLr3h1KPa3U0DGw5rPsPv4cy1F9kf8c0G4OYvP0BCHhDDQ207sp34RZGP7BRVGLB6NQOC/iZ63
kreTgfcKSt7dzsVCTiyLq5kskcmg+to8D+EDkmeycJxeNYBh+vAS0R0+iaFnITXO27e1bTmzQm8L
KIBuFnn0XooQpVLiqgGCtLD4lJC9HetsamAw8kHrSPhwstUid0gVJ0Hq/CSebA/dWTw1jHRF6M/R
08AchO7V5Ev01nazJcA+80ajuPWv/gh8b7BAIxMzmgdgbhZbodIdV0lj3v5YwbSEijCsH3LSGZbo
lfU+1sKXv1V1iazxh2acNOUqm86NmpaR0ydytoxBV5wqTtRa6q+ucy+WyCf61tY11iVbmQVXqfvF
xFWK02BKMRJoGrxcGL88nwNv9OvM/r0GmcVe0wNMx3OZZPG6Sk0vZ069ujJDon0/v+lrrHxnEdml
utgD3kuvH2WhQkkYTObAztSh3fscE39lqObFvLItj8YH2uxuUUOukRg/ojFuWSTC3g61sLs/lcKn
cQZgQ2XXeNC76qWllaFfeGvRPkLcGBH9cSMlftyy1omtiPKscYeQNYFM+RalfSdkW6KrhzQET7og
0cW0vBhiLPlJ2K62iOeHCEMSLTWAL0Wfm/si+UDg8ykvGY4VNFJj0x9ductHTnupmgo5amYul6vu
yem9jsfZbcRv0BTIOQ6LWtHcPglUnZDlLqf0ahqsV4j4P2Kni4Td/86PGnqh9sIAhhvbKOwzcjUJ
wjJ/Z1qIC+OzdzRsi/Vo/u1mA7YR3DVVTBwNytQjq1w45rvhat8bNhPyxL7aQIDawuyNQUZSZGJt
O+Oh2T1IPjOrJbUUUqeFQNGmKTlwQ68VhGg3mswCHlPC/qxwG6M7rWUG0oLWDDCkrvDYbZo+g4JG
hdc6GDH8NTkBRbvqAIs6suNs8O7syVZ/Gdm29TYNriimLIoo5pyR1Nl+1G4RDNlQyWH4etaiaw6U
Z1QpFC3lY5XWw1Rnx8KrAuxApVR/AT4kQregzaZrCX4HdkyMkUASy5r3sjoXX2iVNVwdFYyMJwPK
usS1qA2m3+MoXtkCXqOlv6zb8a/QqsnGHQiB3rv+eCFe3RExMu8lF8SoyXOko06INC9BfYJ4FVKF
MCGgJbheXEnc3vJkNtnNZYHvGpvPybYU4o+IJ1JAw1z+tpA/1fVrJ0GXYM5w2anSyEFLzUsatNHG
c5wPJDuU87ZmSBZpdstWKvwA/evspSfPrJfCd440naThkk24WsQvLcb6EJ7bQ0MbGwGHB7KnU1o/
PV64i+RwN0ns2olg1Y2o7lNr5TBk+n3M/rmcEMxSniodUax1ya6PeCoKhbijXYU3JKYebm+a1fFR
c5vsOTLweRPMzEITlgxoEw9GnxjDGsTcwfJJM+XLQyRlMroilLHR7MVMaUEpELMop4PF/ES6J8vU
tVeR59RhLJvZxXIjFILrwfcKdr7VBxCX8IGel6ZX81jDorfPi/CpAEFWfXqM93Co4SPvvcAeo7EP
KcaHXJUOsmCDVdcUCzggIckEz3VP5OHiVhWcG+EHfQZExGmwymvZbY9i/dS+8snC0jJxPHz/V7wh
huQK6pb38HpqBszLxgIOe/Ll9Pw6OltExbpEPEQfOyhPPtPFYiCX3RRAW3OYHqrbZ+xhZ9ixrkah
oEeYPH9Sxl41dUCY6WJrXoke8npHiQPgUNItniYF0O6KKhd+ty/RoqCiMpiG34ylg2y/2eLkiSRf
CuxzTkS7iw4GD8KVF/iemS48vMGNix7uJaPgDEcBCn28NLqGvYNXcS5m1wnCtTABvQmagRSBE/d0
Twh5DjnYku/IsgtQhALTft53ttmuc0tiHP+JoXe3G4YseMvkpAl4KV6oaSsFy1vbeemJjB0NiI9m
1P+hyKn6ygVehVrdsw6vSNUg5bdL5KNBTE6K0JGB7vjsMqbJ5q+LNJWtiEsVUsavrV5YmFmm1593
Sg8vNPNlkIclmP3ReG5im7mqPQhDpkV4CJplwRQ04yUo45VcvLmz9TzRZkIqaKFC71ud8WJA7NH/
jNe1gHMKx1wQG6d86dzBW0Ny1S4kc5qOVVffHD4wLmlyzSc1dneU8lcD3Zy/xybeS4jOSALnL5Rk
UT60U8hOZFq435qEP8VdxnnCweXUgsPjd9ItqqsGBDvXXSmRN2rK+X4Ljm4cML7xRcyFqsprd8TH
MrnP26ErCUCEwb7vQGRT5J4swFZt/qGwQRXyNx0pfYfdklDq0gVjs9itS7kUZNYD/8cJcgpj6c/D
68Xs72pRGCyPulDJPSDewHbotey/vgTGgu1gbw5Dp4ep1qNx2sme5Y44fqZxw4msFEFoohwbLAdq
razBVw3AVys7FIi2Qqorw4Zs5ws3AOrtK0a0wb32WijdEkJmlPtGHucWSjETuyxf2okJirPhPQ5c
oMN5QBzIU5Ee7eRuxUqicfRkxbc03w0Kfz/jQDLClbee+0RMXJrCwdJHbsw5as2Jk0/9qHQWpPmx
QwF4MVQ195BBSF3vD41aIiuqUxC+GqbqGlabPURfHsCYHh7Y0yIlq7KGUCCJXniJVdIZ8739A9Fw
oDYYj1OyDdI2Ws6xH8OXRjUiJpNjVjVqqGNArW24lQphK/AJCdmt4/66b7Y0MgJfnXyLszCTVnZH
0s+jkVpyT6LqyFOUFspJEG4W1ndQRi5KDylIhD0KaLdKhBwMwIAVAbgChsKayXQrTgKU1/CreJ1w
jX8eF0FNytydQDW2YGeVyExUcMNdnZlWEqi/WvwEEv01mL6t+k65DydhD4YyKixePyMe0bH1Fa0y
3tGz4pG2d9dYDoSTpZrCaUTKcRPjDtnV0YqpORpPlWPSzNh5+71RTAXBF7KVEYre8v4zchEVQilM
JLdl+xoc6dP1H8+aBBVdwFhYa9ciB7Oxr8vCizC9qpyatm+4FwSkjvz/ynrcnAL6UznzzpkO+1Rg
Kk8lIovMtv4ENt5KF8tq8F5qVOjSiJVs6u/ra5FJeEpVaSHmQwFtNdODRgCt9DQlVQjhJC5YT7Bh
uDjzWfr4G9nBsTO8rjZoV9+dJuhLSsV8vjSuMuKPqKZPyM+aRaCKw1/XmMon+krb2gwWrZUC4U37
q3B6akIVQ+tvM+mT863sgKq52WuEQb4d0wE6/oFdbz28AKaTawvXr4FJsRLF0dcFBRy7WFB3SU47
v1TK1mZFijHK6klAOVHgpZnC+wNtQgaMbKuz4t5Empd7Teei/Ioe92d27s7pSxdqn8E7HtX7Be6g
oqyyDgvvSlZhZT9OwFaVBptCT5Gk5MtuKumHroa5TCxgx9fK8gDDz0YBCp9nVn5X1rUG/CTxbkcb
yNZ5/btWJbtT/HPxxT/d8hSNK6wtNrdDGzGmq6l3wz8qVB+gJs1VMdDP8bg2QgtHLFKWkLWgAL9X
sxmUk7uPZXLB7AdqpBwZGf5OYBwjbM4C0yO3gKgXprFH8XJUL9YXmWuzKWKr/cYG8iaZ+zvwe9J7
pKlzo4YvPOxfWKbgyaEDZCfYR4BnEZw88nSkW7Hi+U3rSmsQ57HgRHD2NDyddaBak6UNWQQ8D5FH
mar2+JwmK0pUblOUWXP9557P+mWUwIC6r+2ow4v3HWbl1mYCamWtPPejNkDb9cMYm2G8xcOGWbr4
Fmh/suTouC1DRfEstynk6J4/TIqu/5mv6UVXCK2P7aOd0g1v2uZJ8NV6SbzHzSL46iExhEOlAA/Z
pXZXPJET6UM8esxXanyl5h6s810SqgJ5FlXdcS+EKOVFFJ/T5BqrpfnxGYBNHPERhkv/LKZiGtPx
ftRwbiTBHBVwSmu7NKjN76qIXT9lNqe0D2U4GGebAgGeDAi7oxalREaz1S3aGMNnafA550qb8H8A
juf0PpBb1wz+Wh91PvjkbqPq7A9vpGBdFt89FskV7+Oi6iAevn8TrM6FgVdG5KTp4xDnxa6aiB/t
rpd19hW/FNEYGlkbfOvsH+78LvYY8Ur3o24NM6DwOKRFQCSlyq/nchzKvnw8WhAtrvjXxiipc8Fl
S6cvlZzcp6d8W87gTeELoKhu8X5TYLDwummfvH/g9Wv2KPvY4C3QW48+X4XmO7zitAc8ahUIBohS
Ih1NMaQC6NWMArxoGzP5VftY0JfwUySOxgkAnQguunbb/uBaNc0bG8JIjGA0MPob3iB24RghRB9E
opPzhLxbZ5wmB2WWlU7En8wAUTdenN9S72KcpU76ymxZ8PbGYg3W1xYyeJRS23SUSsRU6aiVt579
OCj1YMtbW416aFQWz0woLoPA7mg4mNi5j8OXM5ffzFxDScXH+3sjQfcvp09hwlq4+KcKLSgaPygk
EYeZq0RQ49sqRyy/kq1o87i7fk/ArHfstUUi/hDopdKrAnJXigBjhIzq6s0SES2UEJcPcXNsUU77
kjP9+agmaHx1Ej2hNwy2fuKyjwxvpftooHUONXkGA/oIYOH49bVjyhGPE1LgbCW1+P1Vdd2TEctp
LhGYzcfp4DHKoeAtrDz1D36yPn6LLXYODrfWePJJKz3WzL9/6X7sE5ebTyHxIs8MvHa8GgEYUQ4M
yrslktH31NWv/OO0KsUyUHEJ4/mSOHt2K7J0V22U6sTFzfrZMW1JEdsNNXsDmrqB7o2QLe/Qxf7m
lMUrG2cTff6VqneU+Ta0LZ+9usYVXR5+Dh90cpJd1osET2YvswTQAkI+PZNQzIVbmJ/KipoYTqNY
WqNz+CvC2wuqA67MGTWOGoF6VqlgX6vtDgV6QQi8Ea/KaliBTczSmOqKXTrTXzrKrvKbmMglFCZy
bCEXypL52V6sSGuyoR/4ej5+kRE2qbBuZgY2G3dFCHdLmUDKPN0iom/yQk7HMEgnG6+jeQWeyngw
Xf+5HkUb4GPrJr1mRH07LyXHx+t0hZEQQbITcOjaIOySqG1eDsrr3GDfoaAH+Q5kycNESSR/+tuo
Kp5N3MJW6JZSCdrL40NZPP6pFaoLD1mv/3AIV3Ktr01Rx4mM49FEPVAtaiUtKXhGtE00V9qju42Q
4wpoMRmvbxgizZ32h95LOYtALnUiBUcWAVIaUMhd17ijAvpGKTCY8kqascUfiCCGWmMbx6prZgXD
cvBIgBmVIVMbvdRr2TZCa+wkwypM8HlOveG/6/wCKIG/n5cu7R5BZ1h4yHwZe+wOsRojjuHDmPre
9unI/TrI3XoiyP1RaLRwKlcxZW6JGva8zyuK+jE/kK7zsHhiInGzCQh1AWmFK0jmHewZYgTXoE1z
ZBXoKOP6R+0MO45+b4cuYmvjLNcdJ97r1wVxLVglbK9g8waBDdNwmmZ9+Un0sNkg5/co9ld77M4F
1X0WpXFI5FnjfzaNGd+AhiLZvDXJ+JaAGB3tZtjE2CCiSniDnMHlGjOU3uzY0+L4vu6Pt8rzIlHW
OTGLphWb1vPjbS2+CKyzranuzMaiNPX+ok2DDcsUeJSWEPqZtU2wdx1DYh4YJXZB7WqrdTUmJTA5
YYIMOjtAO0WXIQN4Z0j4UTDH8MtxTqhnoSruuKK9actqj7RT9E3uxIE57FF9x5aEQfQCu30CitJw
ky7l/iv3HxAmzulcnjyCnOQttten99TGw+0TGetIwwmkj1/TAs9qlaB57X+JMdGI7OC3IvkqMI9R
5BTMhHxOxDxteYlcno91hoveiCwwlkJwGS5Sjcvt4tEC73vBfri4fEB5Ogdi+ffRj9DCzOKY0h+P
S6orrOAi33PhY1Xvmlvjx4cFJjqivb5HORmTwqb0OvWsGn0TTz4YSizhXqhwTGcwcueDQe+qzGsC
tSTFyW9hxmzn2Afi47yz/iHEKh7pDx2eqSRqXB0POkAlId2nK/LHBoeQMX7LO3MNciQ2oi1qzQP0
ZcjlVxFXEvLkOV3EyhZrXnYmeIa+Bw3r4z/L4oRjowVVQXf+Y4ndO16QZlWUJFQXs6td5zAUwwOK
nR22HZo6n2mruDqJF/qmslpBfZX4V5yFQiI3ZxzbNicpC9h0w4k5n4en5p7N4h9KHwoq6DVB8MIo
0G8rcwD5yDoSDZ5BfF4/F/HVO4TYIobCwt5h/V7PlbU0biAcrQ70yA9AZwpCKsAK1g1jUyw6PcsH
oF+9dor+ktI7QYNUepuvjC2PfuZ2OwrEMcnAf7kejs8DHmbNo9z4L+svpXB7E+DDLg3jouSPXBvh
xX3T1dYmUk8Z2eKEiDbli8ISDETmeApR0j3TRju63NhkWakMgsTkMpCiC7eK33y9g62GVehIBXZd
56v0jJvgeVIVb6uYh3lkPj48OOuv40mRAoE+bKed9oasZbpIIk+R/GQ+zxVRCIXOFW2il/X/H99l
kI0mIIdAn/TWvTM6NxCI1UNhnL/AYJTsyS/UJOAiq//MYgAal7291He4hX71WdH0du5SJ7kpEBO1
Mz/++zhIqJdSpmy6/HEduLBd+qoQ2f2c6IWwy3A7TNwttwxejnKdMI84U0mkbeonXyYHGbgFpfgV
4EK2ctCAOz4KEJ7jhe0/MSiB99uDYdvlypsOkhKApn+QEi+aimgFWHgqYgEj5KmVRKF1zjlqxVva
6RCUk10XLbnxd4PtVCWKUK1x15e4A42IIz2FpEA3uqlgHIv2Y/2wUByMFxQOhgKY1j6gl17Q2nbC
FJ9jNV4y9W86GDAkp0ugwXJGVoQV8FFflsvOBO8vJuOGPfTOZ9hG0oJr6iyKuthqlz7uvDPdi8cM
X6LWKjPtCdL+Xv1uMqY1n6C6YbNq8qPrA1OM0pPEReJaJEt0KT0VgHHyt25T2Rht6TRrJk5ViWtQ
+D1j3NshlepmDqo2rxU88+yGLY06YLKH9ORIgWN6t8jJptIoJpRsIczLK//kuzKTEqjBNBEhcRMs
WvBhr0YTIbB3FX4jno5k+iJQzW/TB5nwDT+hoMhoBH1Z+hfjvFRYAV4tD8bN6KK2w8PNXXuCz45j
BxVoe6GdOhLs7qadJYn+GZNYddux6j6je4+bkBeQoBlMGtJzXXhCpASbSdj3LuFR2NXL2UYz1fz/
xLY7y7woM2FBk+R9469lHYvzECmtiJqtYfZ+F/9o6t2CmI0Md95gLu6qLLfeX/pPKc8t1cRab5Q8
K64p0lYriw49HNwAmOJW5xxMgRpcbWUD1E8Ox1meNOFI3axTdsOgbydLpv8BrAdHmJvqSq2kRx7g
uFgIYi4r/byyLEGSg3MCAynULA3lQXrfK08RcLdsMa3dcvsrkzB09qg6E1D4BRoos+812xOpec4c
w+lcv054NLr1/4Iaw1JTh2vilt1iNkyDM7lP5MyPZfdiHjNX+o9QzLfU2a7pIArJ2vFfKJW3vq62
F/zMa3keZdNC/A2eq+yEZpC5bvkGv5uYDigcahUe+Z+hVYSgAvT3rpx28v/I0M0t0t4yVedSEKtC
qJthWXDbMB1N7TjHcbGBf1xU43xmxViavc4ZrLIiQr3q866nzgrbwSW6z7oymreJczDcdtl8WuLk
vCSSYTuqIOcTMaTP5+Qao53fCwOTeMuRmNbTlkEmimfm76s1o1/VECHX+/C5ThwGNhW8EzlBYisB
bI4j6Yh2Xk/pFCAxxsPjPKbwZzS7I3acy3t65+zZb5RIIJJxViu1wtAWpveqG1hXZ7zj1XDDSyEL
YV+PBup7Fs+K7UsmQUKhw5kiPDRiuDBJInZCnmvM6dmS7HSbj51oQhL9ILGYGb/Wf1+27HLoqUaK
cF/hlhOn2StPktWpDxmzWHLzgMCaTY+CKWQTU8PAfG5582X7ADYMcGzbriwP6mC1Ymjd2bOzaMCD
wC2cN5h/hw2NM3MvJ2Im/zIqq9punqvUUY7gjSXLwP8J2vHV6WjBR3u8c9NKUTFk25JSf1WALQ9V
ZL4J1TKcFDt5qIDZNWcQmmGhNbQtC79e/ePP1FvrBpvCyzcUOQiFvxEyXSknJ6HeJzgbAZhDuiua
o+0J/4l9pFvi4c2mmt3ENSxh7sEGbzrv2RqC2073grc85xxT3uohWo29pTSLgGPmiYxRjyFo8ZJe
enNiLqZUsR4HFPxHA0kiakc0fLrdS5qkjzRy7obdoq/UHhWgFhjT4DE7BPYr5ion3rB6hO/YWTD3
CO4otTfA928TetQ6S8p/oqbbDBkaIFL7JxyWDaGJuqglsuOCaiEWmhlmm4R60O41qW7Zh9gGV89e
xivZM0eQEFlWvutvEnDyUFRcvtUMmRDDgE/6zvEPHiMwHf5yE03alQYATIQfV/Z2H4IRAtOsHKT1
J0HkD8KdnyaAFOP6z7ufVx6IQhQJM3hUH7qsbuuYKNKLXbTY5u/XZK2yckcKx1Uk5Q6+dwv5jzAT
CnZFFcUXM46sDvG4lO8skOuRNDJHn4TkQ/gr65Ll+psnQMS7/SQeE8uTKE0rvB9h4uXaxNl/puC+
NXtANGkbuq19Sd37o4zof8wC8Qbj+b2hwaYJsjBYeAZfkfiTAWsv2C7+cmhE2pueqJiSUUJzdGMv
kdzk1937ns1yYy8rs6vHbKhRVT08V8z0a6d7gRfefhAqXjIZaeSSIgpMIKapB5vmhtwOp0WAVOdA
OQ1PhGBz8tQ+SLUyfWGDbGegSQItshJSIl6nWJBRwgMXaBiabOOcH7SmGdvvndW4HFFPx2hqEcwc
Z/7M1Vb1O56Gc9ALXvbVrDR+Ymhu4T1oPfz1tq4wmRNh1v/UhuMsngQKCxED6hicnM47g8hybvsO
OvUSBfLyzK40wDE4gQ2OSjaNwz3hl2r8XRvWPj9Eil3ran7WmNWwLit7NTlzfdJGquBMSXyQIIjY
U3RtZckExOon8Z5QKVtP/h/NbmTvnJ11P92NJoQRcTYsaOao8ykaMAILfJxUhGYSst5/HSt4z53x
G+hUWcLmLnY0++cYVBqqSJRKoPBgZaJHf1q3e2HgDMLD8PdNkTMF/SmEWoj4KSaH606SW+4++lxV
nDTH8AJ6bDVknIsN6Gxcl+SGUJs9cANJA4zvPDXnvMTxmFH3J1p50h/wJoekoPFXGuNGatACF0AO
kwdPss8c0IJKwLMra0ctwXyW+t8/udW/nz64xoDkHyq2GvYRvOntEIwiME2wcDY94MzplckVoQkD
ye5Gf4qK0dLv+fFcsOdiPrnWwsmBd1tWkSrMnqGmeuDB0sIaLlj8XpjpIIZTwhxKqHf0SARFDdDT
AM4ZMDy2HOXbTjPQiDa4qeE62W0UAr6eYJ8/ArxgveHPRGfvYQQPsOuikboX3Vn5NBElvAKU6fdw
I6T2m7xlnHLX14uInb3dN6A7ohmFsMBIH4xx+QFpt63ZQhlT4D2Ys6P4zw67t31jiOFl0Nz47zCN
viu6TOhgDjEKjFDMbpLKUsA5CTakp5RHTUhw/F3dlbsz/U686M/yhzmUsYJ6CzCF/qEZALma6c39
+ZLBnUejgA41KuIMX1gu8k6HZK+hD8+g4iTz0Iz0YroSrhfbuMpzzUxdUUXfox5V3h1QGqD06GLL
2U2E1lsAaH7WiB99AQEjA8VYsrtbA/krvx0kjnrlLHPq37csqS4NQ2CIb+9aYsXd15ftmHpcfAfj
O17h0jEaWg5G+2m4hGDSSOb5WLSEvo6197hB0WqyHFVllH1uw7OcxG/JNnsDAf1BaNC6R+z8pI6M
VZ2PuOqK4yJAGmADwexRJVGTBwcUOzurZlLZTx+IjpvlRRMLZExwRor+xI3IttyMJZaAF2JxOVE0
FWtnQCoZ9cgtBoZXT7y4Y7zzZaLNXjgCwnuZlUXl6YLznJeMz3DcbOMkkboHnli2fQVL6kGzFmJu
uANxC9mldTCrdODlpXg1eflMljYCdd3XE8SuIQ9Ss1YbPo5SNSs0HQB6ZcOnzuSSGKgaV47Y64wV
Z9KA7k40La7fVMsx5VVp53RzNG1BbrKOZ6HOsk1rJfhjqfBpcQa7Uegd228kGq+Kcec6MrnoZ/fx
lJTlSq7pvEK9lxBYqjkJVFpS9zM4VzHoUSO99lKNvF3u7W7KazA7zjiWZZ42RI+EBibh2Jqyheq0
dgW7p/BEr9SMe8/bTswvnepQenCFOe4NResqoqxf1U5nhhCMMZWdmboBX09aCeMN0nTZ4KYSp5D6
YHPNFIOvUYrIRQ36pMUEND2PzDboutez/GUn75fFxAAtYRB1ooucsBV34sehy1EfADqqV2saP4Nx
4JBxLj8cz07/vt5ckh25A4/ewrqPiMyoxCDy+VS28JHexucuRwPYMoAVLp6jFCuPqA87sezAl4Kh
ulB15MkZYxfvP2+yeGvJWvGgYe7DxSJGs6XIc3grLhyrg3G49bro54b0Yc0ocye7C7WY0jZ+jd39
6n17z81BbbYpaEGc1YUQB3TA9ur9NHxwKovE+YkxROzP7r2mvBKvlAxtQ6cZZkuyXT0OQpHBLB6R
oxmRwBDSRpvM32zMnT0Roa4StZAK2cv4cejmzrQEH6nhpaxUbpI9OhTLPQMI8kMP0pr6g6c4fazj
YG7JxVDzwUwBwCHnHa/NOHwgung0r4YZ05RAZvCauJmYFqnJTHF1XuxN7CcUHdLy18NiNCodzIHh
PQ/VTDU/++Jk0drlR98OOdlJbBR8CKYsguCeVtZcUZ+LwFl4mwv4voVriplqkhVT7M3SBrrH9I1q
c+jSOf58k7KwdJuuEIMecGBclS7TXWf1Kl8Kh2PynefMTl5etZCtH8qWzmmwuwyoHoTY3oYeA916
AgYs2GKmX9cfT8AFhhMx+5K1VkkIWL3gPMcuglzQj7imH+JoUDddT3L8Buojy/z/aPyUI95HVvRP
Ld4bwa7vn7JRdRIpgBbX6QRwCvoj6tPxUK0F3wcwInNmdgj1lFLa2FfEzSz5ZBDRTVFMk1sZnyKf
SYMjDMn28bdPp5GxMbW1072bXySxwTLDWUG32fZ3ZaKURqMNtppmK8KiAewuNBU3ViASwSaJMdXC
eP+qZ4WGXhxFTZgX9scWNQblHpir86RpzlO3LDOwDxnpHjGfSnaZIbhzuWnDNSiXaCJiW4cvw2CU
alf2PLc5bLg4Xs91gn1SW4EFkSjiXuB6sbKadM/CKC4sBs9+IFQmgglVgzmnnfIfZODz52BdPNVe
5EvXDTivBVNvXnoQNzDB5cTrZAnW8fBcR+kBcDQTFpoEiC4iGc7Kkkl6IGKU8QgJot0RjIaP2dxl
uwj+x62K3Z8Vq+LEGaGeKb4+ojA5DYLywu+FNop1k+vfBE6zOS36HuomLhdwBnB6MtO4UKrK7EGe
qlTd0R2bbAEf/fhWDMpjY60sr+iiJ7qGLLxm4A5r0SUKv1S2FtwVzBnr484xvEfPLyb7r8wc1Zio
TfdUVf2dYS+HWb8rWiteQIFC5PDLAR7+8QAs5xR4heWGiqQPpXtnmVY+ROIQUvpx8zLQUmhpttfe
Z7WBMivEmIkg2jYoF4txEMU3gV3UEWt1uW+l+mVsqdGKuw5QrZ8Mg8YSdH2eNPTqTKz1jSmbngJ6
IAKE51vdDR/nN9D6jPYFhASHTZK5+8fSylHTtiWZqn9/EDctOfrEfbBtj5toQqUOtukOl8i3MF/r
KW79azxsdbzvxklrtx/kKg3Uc0kpQZ2lhK1bNIeAUgbYR0g1jPrWTxKqEzsZ5VCimfU1HwjSi4un
h1w2vMGkwOAyVy0RphepDAp5FtpxjEY9M1PN6CKqRfC1uh7fcib00HsEdqEbRb5xJAeUzHKA26eF
H4LIrUdWzb2BSZRZ13pkQVPPfoNs53ftiXYQgGYt8mjrrXNe9H3vBq0ljh2cbRANyXRPO+NIckcX
J5J7EWu7QtMEtQftZ8GmHku2Q0iVZUOVV+s6f8lfeW3cthAFvGkY2oJgbpfZfpjx6R84cIo6JLRl
FXfUW13/CV604Vsy5oSymHJK433nPa3wAeeHwqIF/lXwcB9yJDPTCeN2ng6UEd1IgaVIrzlO49CE
eR2XBDaGfgfRWyRhWm6ceQ+Wa98otgvGg59Tp2O61/p56sHOq5dFEYoxFBDY5CbiW3qpunlje+TT
TnMBtCrLs36r82NQlaPRqG0ACfUBr55cO1Cu81PIqo/vw24ut6DTAc/JTT4o60Rp9IJY7NZYH1dY
jFFXCqKF/fSi+I23NwA7DXrvuoCt/m2r7nY+RcaFcZDOIV7o8ctUnDaWuCTpEWEadrlQRh+9iFA6
gN7UqPrvBcKOVlD+otsBK4+kV4sbClQ2g6tEc5dZvimNFupLRJ1a71Pc9eJ+ShActplhLM4LMypj
Bm15gjE5QOEPyHd8PrI9dJzip0RQMs7yWLRJxzecgSZq0G++5RClSG7/x5D2omQFJh/gd/5ZelVP
1PLXohgvNUHQ/6iDmIB6HJcgnEF8360oqjbwoxo11W4FZ8ha9GbUwBgx8DoYCclCTeieUTJMGy28
T+op8cyLkge9ES2vPdWkQ4LrEe/zDN1IqBE43mx+9zrp8lBGQeX0ZUv3q2cH8dHS3/XgEQwDCAP0
CfIOicf4TzlHhHaCqc1ouSIQ+DoRoDK8rTpcAA1t5ptuyIh+KKAgwdoxhXssphvBivEUqiwkslRX
NvG+L2Fx11VWhVXztIh3A8NNvXTm6aIM4gv3gyMAczrkgvLhheQ9VAMMwmuzXdhkVj0ceQ6d0z+0
eKofGwL69Iluyf/YBxoXasjx6OxiiLeZRwrBe1dzbhfbpmvSUrDw2Xrof5HKdxvRnXeeX9jJbszd
QYhjW9n0RbJ4eCe4eD2xS69eOvGiBxu/m5McdaIgSctXP47X2fcy0XW+RL1fnpcSyDvJz8zOK4LL
DUp/ZBLQszgExLfZPALPP41nyUj3+FJVHv9TlP3ETk3c/vazzW2o/p4k+TyZfSy0KzDoAEmqyOQd
cnSiTA5gPwiX48rzk0qOQdC9SMx9uHdONfIJzG/Qe45ZUIRk261KMbRrTktZ24DxxlwE9sQsKcMa
0+xunLikokm7GPms1GcoCkPRhvsurqAKJbW2GXcxdPbvybW57wUaEGKs+St/3yMhbIs3EmdWDg2m
Lw5xTPTBN9knjHknkaUtNb4M3uPZmNdv/q8+v/8sXfokaSOCoRF5t7RXgPrPaj2YWG4hOrBaaFvJ
zASLYOQAUXmcnGy4UTk3jcIZYesIY0xEgWOTIqUKTI9eSo6Xdx6O0S6nuUHTYkmtKkmQN32km2k4
yEnaAzxrR5mcWKpIoNp/vd+ecQOnirPKrEYfzJLrE1VozY0J64XS7pq4mtKtBpyyyUb8daV3Iuv+
qjUHv97Uih8ZyTzE3H9p34bMfjx82XytQOq7vaxetzymttscPGhWh3A//ojYlh2ln5eabyU19wIb
PK1jGhcnO8G1EPx4QYeLVSLX4glf/doFGbXlifFqE8zlKDJ/EChzORFDYp8izVEQONLYc1Sr5+wm
yr2uCGYBn9IKkC+EqJCrZ7p0r/kb4qIWujxjCwtmMy4TbmenwDn89no0neQgRmd1Nj+aHYtb5K/m
Ywf3jFx7mQ5+zZfdlowu9oPcyjEDq/NR2a8WaCEitE42qE/QG1pO3vBKUcuGAQLzziT3Q/VgGgWV
AAMG9cxDWwMaVpmeQe3XlltukUrqZ2v4BaEIy/3ug8p0tBNjljDPx6/gRA7T+gLWv7FzlJEtbZUF
IcXy2gT1YQMn50yBQq3iul18zVQIh0wFybx9VclUY57mfiT4cR+uiPIi31kz2e+l+ZgABNMeFL6B
V93hWnAZPmAF9IWkgjlVjKiBrRQonYyEbPkv/2AyTmhvZDZpvF/Qx/JMw/w2TxkfpZrpvFZxGo83
Fr9x7rPlDpyhawsd5b+YTmZBFTsl+r4+wBZlX/PoTsXddlJ1iptIdRnFGIthkMbLFtaEaRzfeSZo
HuZXqu0JoS5TLPBVnhK1IqpB6GsGcGFI0qSFBp2xekctn12irTlW6V5XMKcRotiIq7wf5FKuUIjr
vbtqhTNo2yRPuIKko2WHU+eFOCyOGN7zdxRebW+0KuXbfTMDaE24y9DOxZ/wehCMzcHHjU5Vpkap
Jx03wDZby0RZCyGMrgtboF4uUBnX/vT499Spox/gCyfeDY5NZiMYfuMZ6kkzBQBus0aKUpg5bNqp
CaZ9wea+6Jo8FUSigvQkLGFgnLtA3/NvYhWbTt18b0BFXzDAmkEeG+50JXWMA+Edanp2xtMOLU9Z
lqu46GP47gdHToIBtbMkd/aDgs1gb4xouY6yKX/kYJuji5PGqIeDlYjfQEubGRTGUMe1Kxa5RFFN
bQr3l/0e7rt/2kohD/wxi8WosTBc5fvEbH5ZfG76bf7vAaTUYomUYcqF12wEdVmaFVOLDozvr+FK
DnqO8G9xnmMwjTMEBMC9FcPTr1U3/R6EEMV7QunOmbeFEcPi4rqpasUIFCLe5I5QfLWfCkUVA6rV
oorLb8rYdI9pHmUYyw6ESkRS6EtWa76UgKcn7lmwb6HSJDzx3U1C9LMC0HfW6WPoM0DcUsOVPS3a
k9VGkbsx7WV2x12yu7H+WyHc/K/ye2KZ2fVGbsLiFr3jDOfTKCCDxlEJzfBq1XDgzJJxOqDitPPw
tli3Ip7n9pDX83pUnjcJIXK38Uu39f4sykU77A0A/N5cCXGIQCb4ZufWwwaP6Xe8onmUSNmodCJD
GUaOKDCRbF+9VZGf5ofZDJEQKuicRo1Qpp+I8ZM9kDdBms8gQg2qYnZxV6tIwn5FUMzCOGfUMVOt
EXtyriO/TzI0jwZU4VG3sWTIcq5ZndUk8lmdi2DlOjkBz+MN7mHicAk7mNjUqyM+4mRjWdHC05If
Pt6vDb92EpaAPNWverxhSbfybGEkvtqnNcMFq25CGmFhFJFfKeJxAHYTjTmTSXszaG7VEDhZd8lI
mkm+46WzhWbstrrx1cShyxzs+jyaozabQHJ0nfe3/NK19O+wJE/0qeNm/5f8pd7okvY1G3//jdGj
COi3bTWemJx+sIUBr3b6pI2dJ0ivahrTYYS7WSKAoI4puN2aHT7zpSp9Edn8DOUk/HCfg4awmobV
STvhZqP8uuJWbHFUIarQxLmLMae9LnpgOEMX5NIynngopydYgLOmVGmWcsYpxonSTJwHNlOTYmqd
RfYO1FfLoWeIt5Gt2md0qmX2U8kJojx0+xAyDRDho+jWR72sYPhRMAV+ia2DphltxIVqbHbJQvBj
N8O5Aoaqa9u0VEu7ylwmg6wpoSJDlnRI6tqx2w4NWNarloBZLCTZG2wUQ+Z4VTdQ6VzcqJ4OnQOW
InBMI2NhGntzVkzWbx6e0qCoPg0cxt8wNVe5PhG/uEfYoY6ST67NGXHkUaJnkILLb7oAPTwrkF3n
GQmOm+OPgcvkHcMagr4KsXT7t3lur10EO8TWM0hEcroj1jCDbezK4LOXcgEkTV0jdmirCe+xFn3x
KMvsZn1qe2rjsqcqsEm8gGuXWyE3SvnqmvVKXyII+4Gh/+adFPPUf/L8i8RrF2L8GTnQ44g3WsT5
TZUtYfoG67GlggYUZGWE12Pvp9emqCuOUNjhRtMgAfwHN4biJNSP3YU8b5RehIsddWgpyaKuww/s
tzwNEKDuTSzTEqurUs6nxe/Rgt7vQJ+SEIMYv2QV6wd9Kb+pfANBb3LvsWiiGNPND5CkPp1aBVCX
w+WzXeDtjGdOsBwoW5uSv0/zs0snWG15S7uZ0iyOj+aB0lZXyu4HXAm2oHqAnnfuThbUqk2hvQ1b
r199bic7pUkOgqUsUdnbtNfOSlGv5x9e/D0hbBGf+UO6xwOvWmmeo5C3ca0a02SqxNbsCUIZk6kc
lVwRkJm1xIrrvYliCDiYd0SZyeYI/j2/D0YiQfLNwlHmpjbKtTztAh13IJMiKxM5hEQQv1YqQwyS
AAw1tzdxSJY0PGtSFogt1shyx9PCz7RAIUSCTFCGJJ9jrCZKRxKM0Bnl8eFApPkBd/e7AVlpxPz+
VVrZ8E/V6aiWiDZ4hQ8fPJoXhWs2rw035TUycjhUm73sHgwCj8qq8flgQYs0fxWxIFjJ8GuU1wbV
+aljd+CyqFB5nteGjbZooUmwshOYsTZn4IkPprF54f8PF4/j71PH/o72mLPD+dGPAwLoZ404HD/9
74lauTNeRTPRtQaRgD+vCQw1nt2a9ul92D0vohhzrhET7+xrxmKAWsHUbpLi/fPlOjLkdBy5TJld
AlIVHK54A5YbmGeKlHYPCrG8URIVN04BwsGIUtKwHyQLRIKHMTKhj6y3sDW+vse84Ox8zW65Z/t2
iz3BA7oX6wsclbrIHU1n44tR+clGmySpAcn41yTvayvqGmoyFoXWslO0+otDmUHSLddA/cwZT9M4
J9KQIKsdycwbzzAkmVOfM3KSAiALIf9lIPiO2DsH3Aj++HSoUbuoMeY7BGUg9DD9SsOgNFXMQie6
k2DfHJGyNdOuzUUVGxfj2MMaNaa+aSKZrvGxVE2ZUig7kju9zBP5xgdZ9R4IZclSOAxNT/yco3tE
nYVKddz6OiSxFNn1PO4FmX08uhxKmlM6dv3/hbC7kHZIiM24w+YT7hTdnBcUDt8KZHouGX6IWO5H
6VKP9eyzj+ualTgrI+vwNe+ihh3gIz+DS2CeJL6J9AYbOI/8yJlfr1XYLlRlEg2U+tFxORQv5+6o
vljTiihVr4A8D/D4B/b/Pm6xX47+JlHAN/nacJLFhbY7jtXvOfQ0DCEEZpqxwZUxV6WL1UIWjUXH
dSBhQEMGKnCrDszJGeX6AHwW95gg+fspT2w8dIuqQUb4aLYh6ygFbY36mnGK1tlRogpJjRxNjn4d
7rH7uqdylzxvIzxmwz6wy8KACmQguoU3Vq4e7e1AmSkSTSKpYTZouh9QaG9MtxA0lJ8LL734ZB7+
rUtK6qyCMsHrwknD6DO/Tk0ghzLmdTBV+BgzT3EH2vnhiCCYCFf8LBHlWwbOooZ4AQyiqnuNTYwn
9iEAHJ6fKYejoT9LgVXBXxtGIBWvpS0E2vtyjnzN9ANmJ3BimoQ3WFQn7EDq7W7aD6j7TRhiYYU5
WSP5U0fZCpRdflP4XiSwEetmGIFsS4+ucqHgY1HzDrpbd163R80MDDzOL4UyqoX2ApXLT5AWGHZh
Tlq8XD354bWHE+h8fJTacdyiHAboYeAufVuwO4+qb7jsRq1KqhBX95+R/7cUsw8NgC7PCbY9pcLD
qoRVIrQc4flGbwezVjSTTU9U3+I2ZgY2SenRK36rknf3swy5+FrNjG/6PJLqpXGq0vIRQEjrhVAg
C+XD8Lr8qdqlsuU7Xb+HSIoCEv8MYwpXtBE+hJ4hd8WqhyZsACgmFUC+xrcyzoUhwJo1taf/GRY7
ebxZOvWPPIJcE0jxP2aP5pUgA41hmz6Fs0ZMUtqjv+e0cN3WejxmaWwBhsgLUXI+9CNO/bd3w7Ws
zAj5+G2iTZZXBSt8BB3aH2J/E4Jb6xDW2T4zCpgLfnIAOSXSJxtp22P6Hi31Se0E9O91yiM1zzwI
kL0K5ciBoyAvM8qGDDtzRAzewrS9IOd6OLq29jI6eC1uEDgRrTaNP23R62/wifbKkHvP98+QLdOq
GoVWRSaIPo0lpcYF/710I33+RO2M2yn/h+vFNMsmoEOsP664+JSRtROfd0G6Tr3UOP5V9pyE6IRc
Lmw6xql+dP/HVFz3HKzxcLFCgAkKTjgrExemzDucvNMH7qAIfH1GThEtc6omkQWxUhdX50vMEr3g
MoSVloYWX006VgDVyOFHfToyeuj37gUYYSxrWLc8I/t7nzoixWLI8RHrjUMTcuq0FOtXZ3qn4zB0
JNWLx51nJOeti081bpr1NmEGkRfclykWyU+UW49Xi8s6Colr78J6zv7jNymO3VkCqnc4WJPuL1kE
pvESaVeLHfuY8HK005QnnZTzSgbwsHuDUzDE38/rMf/sOuBewZBAFxCTyY3NxNxDByOx58FJdjsH
b6UcZz6IBpbmEyNEvH5qmM4Swv/YsNG9mDkh1hIqUzj+iQG6PCe40tGKPdvGYJiwcjxMjiLD2ZuB
ht0yd164L8gzJkLrlavUYI50aXNG0J3ayqsbciyFGX4WHD44bnjfe3W35x+38QeUgSsbYP3lMNnQ
EpXW1pkoVRzR+xmJKo2hQBULSRzogdrawa4trxUc296Ajo0Jx+8iQ+kbNmGgzWHUvnHVOe+2Skhm
pRKaxiYg2JbqC7ztW3NDrkg8yy72dtsiviNz5KJDyQJM6Rbk2kOAjPLyl1L6bAXPlFKila0xU1Q0
3WLBKU4pKGWjMCp68oWoQrDkI2htfWfE5NUganbq25KDLJq/dLCjtacvAYkkD0TFx11BeMe8l1tu
v5UhtEomm1By+dztNj4kOduT5eOMMH8Yzyhw+zz6CEV3ISJvA8TfONQ1qoB4gKKabGYuTSsV/YSb
YiXgFPVifF2OPKd9Yk9j9LPW9diTw337CnkN1NpWiq1YSRB9QoCJ6fu9AzyPDqzmeF93P3XREJ/M
1YS7576Ls2rgfFhUSNsYT8uneInOMoL4xetWgSiBAPzPrDKraO0fNAKrvVQ/+3EM109TSvwaGZPt
Lqtmr148yMPS9NVaR30bOAIYHMurYDapL0OHRhStBIFQRK5X96T9WAunJUbacMubU9dK2D9KKt5A
DdE2O4R10QH63TESjhaowXeqhnftx5QvAQWDj0ocSH2ganbq3SNajORd6PC0ffvMX+MvVh0X0PJA
fy62cSti9s87xl/MZxJu5+2bWdq68sSMPS3lEELjkLAIdsdeHz708tv1TG6+C038DS89fHBuowVL
oF9l91Ry7arDBhKC4yCSbCh4Hu9tEuu3AuW8DHGvI5VNhIk+B5GACfhPzvDft7epCFy/t+FLyDdV
t/n/qMrcAzpQfd2oWxmEZI3sfOJ7abdPDnTpMnjq0CW+J2BrUKC0GDIbeaE1A8iQ2iCxnjR0mQav
UrpF29JgoBUGackPZNKhnQ2/htLwbOgnRcgAnK41fNydR+RG9sXy2B/+NVBC1RXzADOMDU667fd1
CmxvY83P1RM5z+TwGqR4B/0LL3nA0neNTIYti1qwRu83RRCMlCGx1+JGtqWmnhqxpfJVGH0qAoII
jQ79eDl1s/SVr17ic++AXGAATO+EHNRz+Ud+SuyqnnZ+CpPmPm8VCFHw0LTa7xoHBSOt4Lz9Yd+M
CxCkHtFlOkMTtIBQUXqZTLzpGg9MYM1DPQ8vVepw4uAVg8IxYPzhP9+6+BsUJBIuPxQPF9mS4Toa
I2cn1q+se5ZywogigNr3PrJnMNnwNOMNgRgNLbmLKmq5RhFU5MM5IlretROrf91J57RFmzLUPbnz
exbKAlFYTPdp4NAAohQ8n1ok2UjWWgMuWL94FTacs0OKbPrS0p4A+n24gZt1icL67Q7hfmcfnL6z
ClhcDaw/ApTsaoZjaXIDlTDGCqIB/DQp10r9GZGo4t+GCxhL0/6aUGCulJrK7aYbMN+y+l+mmVQj
9EoYjKvEYj8puwarEuUBnxDCztqzdT0342i+R1l8uFVD723lRBwVasrxniArP4ExRpGTjlUdsPZ/
qoFelqztSD6etfR5fNRoYCR7K9/S2r0tEjBxDXSNbFCsYgG6Z92iZD7+cEcMQGTaEJHWOfpxhc80
dpqiHex8dtfUu93pkjjhzu3ci761OU/0GrZGFSXcb0etN8IFtTg5DbgqE6zahqsabH/e4fPxKuf1
Uli1ocZxIVdzeqbDmd+FE69XpCdCviPwme0LbYluP8em9uX/YpR/avWNP2pqRxRlSAsjayAQjMsp
rp8nIZoKKoorX9/Z4F9mCqrikeLp2pPGPDutacqRbCADH/luy/sfF3dDBxwuPNNRYJEI5ssQt5Ba
/zFnx/Atg2gYY7+90S96mtY4S7/Uhw/C3n2KLQrIP55HHuCzAP9OFEIQ/25UdsbKJCup5wc1PK+o
IfV0mMpZPJJsgNyIp77rLtYoag8rZlyh0PZ22pb00Ex7Z+0JgQkpH2mkaYGJufsqTCrCJV2NyGsQ
vpZginFQUavbdTi4YmU3x9rdkA7F+n7THNzo9wwoElVHtvb8glHoDh5XXbiP8N28iOvuEGvu0fgi
bFnqqBIkMsD9+74eNwBDyxXFKIXe/U42Tvy0JidVindMiUTwHDz9lfx0rEEx4g5iHaXWOzLIUstv
k8LDzquh0XPtgW4P3th/uU5kc/4ZTY68oeItwH9xxCBsmCY21f42gS6OVMnXsxyU/J672vZg7F4H
4IhW1CujfGabJw63PtuA2LP2i4KaFiFyWoRrdCjtraOOAZehpsujsXYcpYrbBj0D7hNGx2DRW8/C
hMz8gNRNXZyOZa7YTAtkHjaXJT2aJyKeVsOzTQMiNYMIDTi5O50FaQLfRENS4QMZjiFdx1B4RPv5
57dNK5BF4X5dpKbAiL+6qh/ErUrVOdzuZ6VDgmyvSvr9RWdE3yW7GU1WHDCTIu9aOmOnRfIsiWrz
PyNMVv8d53I2CuwVNDrap5GtKCKkQyGaT9qqlJ1GE9BfGxZU7rETX50jHq8rACKa+q2iLocFvn3p
AdP8Svt/bSzSjoVL9iG+5HPEMUZRuF3ixGDBlTeMrUS3ABHLfihA66eyEDq6Idg3dl9nOuFb9r89
za3cKIT86MrlcXh1xelLCaqDAsEMZ0WeMGG3kHp7tZb9iIDRV5QL40cHGLWWY81D4HFOibUxCxFJ
rIG7u3qpB4F9/i928q1w7bsrgFPrs5K8R6DS3U5AgQYiAT2yjKRKAl2reESOoEBAe24EirzJMCPj
K0r0bjbf5oIX46SFHUtHsHH2sN77Oj1quEzYUeeZMMxb/PvNLpmnaXRPmm3F2RyCpsvKkvtcTXAh
w0HbGt9zzqFreRfycxF7m37HpsAJkU6DeeKSgYTjoGIP+RW90Ee2MARI/J5AjgdrFQ/hL5MHab9X
i95neO6XSSKW036YY0/12/TuY3Pr5pB7BVq3vpqq5jUDNbMCqmsjtN4kfyfrw2IfEIXTgBFPaZ/5
NGoETUERJszHnDkAWY3Yos6ePVB3hX3Zrhm0F2hFPYIZ/DGdCPws86NiezXca/0GzaIsqOxDSiup
GpQTJeVVrPm69Za1zkNhoUfT5q26bxyt7oZiSvBJmnljsrlHMFS9940W79hnKF51y7Ac6KiU4Ap5
iWh+O3tEfZdUgWIA/iWi7mzxVPMus7vKKRTO55qT9d+3MzHmlHhRCStiByOcP8NwgC9aHH2uqbYz
n/o6hz9NpUAt4ZsBs+QajyuktVCB6J2QWn1VLKZAnWR7tE6cQmL6PyoFfpKh3EpGVZQy64TK8mTz
nePQkHMdtndYz7+sfHqbyU69FwNAYaHG5kvWo9nYK9jBTGFJDb5QZx7aeLiohdgtKUPlnRuU13y/
8JmlDvwlG3HMG1QDMVjpZciEZrmTmTrhdptBw9utZVmAgEwq2VYgi0Iza+cNMzxwRPgJCOTvnY9w
ilCy3HkI7g19n6y0+iQZxII65ETILeLtaTc3Mmuweoql4fJZV2AEhlr2OXog1Zx4AMfeJBWYqQ92
u9u9fksAihgikISIrPjAVK1QRk0tiprOl0c3BxypUf8jIuJdX8Chiijv2tSP6m+5OJpz/5qFBO3m
MFhFphIjAs+BrRj1QFfi1h2AFk2wZDJk5n9yZPciF4QqPfCeMKAwNSr6Okbhxc+Z07O8EVEo6hjT
wTXdw3KMPI75gEzZqRrupd8JIQJ4ApzJ32meEHz0IDVDdz8kuIWpSFydqcIkDqSuubD7nuR1QWka
bgJnPkmgBGYJvNmqYzcvUGGS4vTzipL1EvsQBJ/6HH20YRNSTetLiKEQr2zEVCHrv5VZPvubvF70
Hdio2I5nJTdzQAqzQfkhCfB6G4fTyIttVmeDZ1wis5A0gc3WPTuHDnOZcwt6ftp9WHI7jhGdSl36
7+JQKHQcBpOwgKpbL09lZZ8pnk45E2x/C47I4koUDRAYKhQmzldu0n72lZnrAMjTyKuoUx+/l06p
qKNIRXeBdAZdP+Ss7xTXGhnxG4yRgRcWZmdr+IaCle9QR9U4wUmL3D5rwdyZjogWDUk43nhECF02
+bGYCcA11YP1huhIy4POq8Jsp/iAszvIhNaPcPtjZizfOnnoBv87ycmLFu0UFwPSrikO9rnFA66k
waIggkhu8pQZYXFE61ME/Matn/YMPby79f3burB4aQwRNI0XIvLeKPk+aeOBqfR7q6/rJyYLu3rr
1eb+TCMQL0l88wcx4bInSOGdJeCSqiqED6lgX1Mi9EzW81agYR1NQ6RpsRMCsRQICeIbCANwAF5Y
WiSxcsm1LtR0dKrEIsDXhHr1+hJhoBiLvKlQhEkP+Q5xIISUQuaL8rFG3VQUrIUs/1HALs+9HV8j
0Qsrpt7bBsw3ILp9AGWMHkcGo4UoVeZPbDgCPGIernji3sIWX99pR7x70l5LYGzAeSZw6PGD/RZY
POkhxxCCtQATbXlfLdQ+UQJl3Z8aMbxtIMUkqQRFuRIG0J9+RqSJIV91/pZcufBQPDvX3IoNGPtb
EBMsALDbYPMhY/gD6PzCJE1LQG6llqunzkOgldbEV2Dv4xwZAbU93BLUKJ5xx6rTPLcqx0JLmWdN
fQTZmMKVPh7r6NzU5i1B9D56ZiDXbhWHA2P0ptQWAD397rTuriJBuxuuNh4FWtHR85bYM5yL7u+9
WGUwo3qlcYCY7ETYiFKmfDUtZ7BamtpTFiCYlLiHZlS/5f7jzAITWtKiG9+p3W69yO6VdRUIoPuY
b+X7Foz94SNADxcQW6u9BRdGKTOafWrvvassa77WZ1nbhOtMMxQtBs9KTTuNQz3VEwbEb98t7E2K
AJw49Qv4NPfnmwdG2h0TfoSWMN+kCKB82peDv3a6vXCjVwMhl189QtO9H056CDCpnUM1rW7T5RTU
CQ6MjE1NmiqNSHdf4mq/uzIMgBRVb8sYZHezSdfKKQvyDA4+hvq91lj1lPA/OEtCNuRYrZnAbf1R
mbhIBZsZQevoXuqx+sNuT2MDMmyEXZgD/USl3JZDGYZcfN89/zUMnQilZeH/t3Xb4AYQh6qtykIZ
n8SQVy+ePph60bAVHLhw5odfYf/FrxHT/azApJfXHNG/kzhzu80v9ZxEFwG30fQ1HzD6Rqjtw4R/
eNs5sld9y41livvdi8W1MYIIJ7KDtMVE3PA/Ta2zLcYLmPiv6PZ70z4ByAfGEpStqJbNLhmk6SsG
Bss+vUq3McfpzAkVivBumKhqfakRlFtpT5Z3lvTZVwoUXbPYjZbmuCPf2+qORp6Rogk3+aQz7ASF
BDgkOfJeSjBphYbvw/QqvoWawmiWHksSxhu5UY53zCG5q7l00PNrXBZIwipNWkncUouyr+ofJthL
EO4XolEH4D1Wk8WoLcmLL5mhF+lI2JMoJOc9CJ2Nr8eQPfGY3XF+3FBp+HDi3V4w1slVlcEUSIQd
dhP/XKiyfx+hjr9A2yhLfy8r/4nO5cP40XSa40J/0U+wuxLR5LYXrlHxL/+xRACrxdAmvMTq+Rhm
M1LEPb3sIBDFlHilV4I41LKY7QluAaSGWn1UxWbCJvCsEeRZ1xMv/DrSOw/ZZUrfmXCrogNJwqvt
e0NQExVr53cZVrncNJ/kqaQ/wUXKwIh9eA/2KgUUmmP2YFz9kKQAS4S/X9ysLdlsYJfrVLvIsDtJ
BE2ksDaWngQnkIoW2LzFItnHHvmPkV8byeKcIdfy6UTDQLS4uMVJTYkv4MJL+TQrbUHq+Sw3CqFJ
eqOmpoU8Yt+0dpw3/gpsrSftVUmAMFH1Rd2axrrGzn8NOtMlcN6RDBkHtw1uYqCEGslb6wotZIXS
cvqkNoqopqdKGCvBqtl6DerCtBpQfntvw5pyunMkIFyVSBi1m26v8Vgzlly7HwfkQHw24vTFxH+j
HbR500OxM5Yo/QHpt1sQCg6uzwBIenLEOVgdK4fENZZnT4At+1sYmLauwTd+Di6XPbBFDpcT3bEi
BrS6thqM+UUut4Mh6SvNjLzoWwrG2Nw+x5LgB8yITAqcMEpBP85+3xnl6ewjhn28QuP9vNymA1s6
nKweLribkxmiuOFF4VsvgHBkfkMHyDECdjhCUmSpv5hsdv0EXOjPNdYOn8ZSxuYwDc2xOS43ExdT
Ugej4WP97Bozd1G/gVz/9v0jKWTixZ/7JtLRr8UIRxpdLToc3stIMruTk73YFKUPcqhOkyMR5qe7
uGDrhszkCWU3tODX/AmF6pGJY+6yJdSmlPFYZoysqjjpWvTWpvGkiszeHXeLaHmEs44F2sTL0+o4
I4bMqHCfjUEhz7gbP9cwLjzNg17bT1abCwRQ1/ardPQFBq/TwJhlrufxZJQ42Z/RPC1qgjhq5OP3
51mo9mKEg5XART8jqKN2RfmqYVev8TInXxHHcwQIGPlvJc/0YCwKzWkaOHXgset5ozbjrY9C+gYN
+xnd8XALoDTA/JvB/JyBBttSHHZKpohrQqbLdxmd7ZpMexzgeemuKcKZkwHb6/EgntSBA66jNbEQ
rQ4R448P6TuAAexvnBCkEGeXz0eE16nkDA7GF8qoyWOzma5J3BAcW4ImUOrUQyfZPBpyYS1ZA/A4
N73lYZjTjLqj6n5C18mHLr74ydMf7UWsWbeu4X+LIfbUsxOBnv/uYhgGEo8GzU3Cs0ZgU5EKtohZ
9ah0R9SSrPk9GC8/93T8mvvVWJ2tI0Jhmgo0nI9lMk8ukXpZAky26HusnVh8hxm2u5vjLC1EVXo+
hIeVg2Kg+HWFkmHbAsWZhUrMj0mjZ/z2WQdDKET+fioppOHS5mjclMWIRvy7dvIwx2Ib3q2Nly4y
c+Zd/bzS2khr4eTFVadNRYjMtQ6aFReK7P3zC9Dd2kNUCp8IjjpC4lerxVuPvwwr1vjhRKkiCJ6w
WKBaq2QEnWpwPmwaFJrHetAlASsD6ZbcFlgXsaEwCGEOqhqHC/4VKkdbgmXwihcl7zLJAXt/46Qd
LPQBhLLtBRTvJw3bIzuvVYvivyn4DagAEmCovySC5Qy/WuWdSPH2hbZbqiRL95KIpCJXBqUW+eQx
MpMevKQ6DDrWrUfbU+8kM1+wy5JFzbBp979CrQtxg/lrVAn/T2/5d3G92HLGT6V0PYhjNSwb3w1b
6q2dEAl4qrqtSHBcg/0MWbzYBH5cLhljcUhoU3ETlOG4Hpp+ELEJtu2P3NZTr7/0TXw3lyG5/sGD
EGfyntMkuPDVqGE5wl1KDviWQnqKZKh3BK/CTmFSjpHAh3p3ia0Qdg2co1/txE8tvrNFAcp+2Zsb
LtL/IumivXJCyZLvwkS9uzZItTeM0rpn68PQoiui0B3pEz60+crciqGKjApC3uOqmgMrHXsJKSbo
l4V6GzEg2LvoXk7kRieiQzvQGiPH7GKZuKOjkUCK4nMoend3AgQID15SAXnLFx4QKQ0ht3eFOgU4
rA9PQtNrwJH94gZaKcpIhvrw1wV9n4qkn3cm5VciFHUXDatXm5Su8Ft4NZfGVCxOIXivVxBjyNHE
VxDOTHcLcPfUTcDVXaYYGEnDW81oyqklahD7Nyj0QpoWRPnPq/CgH6gZxcYvTuDLOe/N9MFs6/0L
wdA5+YIyAR4g2wey52oOIcB9QzfcNXpUZx8pvQy2eV66I1tLnizfO1RSXqjUN1AYEj46E5eW8nVc
lq9KGb/HXxV1DdgQJp+WhgpF7KJE4zKrDu78B9SDLjHh9tQ/t1njKyx7cCOJBupQpeAVZ+ecN7Wi
3CqMUTP3RMsIuhZZDdXY0OSBIb6i1hNXGjxM5hRRsGGE7tnmXrAMiV0iiCUK2faIAO8xA+e2Lr5U
kd22rHeNqP6VuHaZdaF8tGqaQe6zH+3P+ZK0GvbyDSl6IvoXtbIKw1Xyb7vZ1WkXRr/+tt2MBvyf
EnlXP223csBu1aDn6pPFILUwx/PCfBNe5SILWrW3JdIvxxH9XMgEm/XJgpDk4RcTd9SwrDULDT/i
uvcYaine0Gw+9r+0LGGtoDeDKoAVNw9YrEKGbICSZ5RG6SbWCR3IYCSbJufd/VWez+TnkxiJqBQN
yO29H2oKFXFCdyyyOvtYmhoqlql/o901gH+QChtft/NtBIEU72a1H6ouFW6YKuAxZsv11db12MQo
naQRKW55/1d855I7i0iy5DrFQFRAv3XeQWac3MKgndhm5qNgoNPtZLjNjf14+BQhUs6eI0Oe9Rqy
sy/g+jRz/sLaIxHZ/injtTuNwK/CjHdbQJgWr4hwROo751kg97BwYxGA7jvsqCqm0s8yi59XQ83D
PNSWYlRa3slwDNwWP6XyXHduMHGZhEjytF0/d23qR20qgg4IYFdp3v8nl16vECbKaulCc8TKqJqy
ZPfBK8zFwEczUXx95etaH/LyFwwwZv7119ZdTb02lq94FUSQNgpDDj3wSNHPlI2AypqARVgICwia
YjyEEJbU4h+tdtxLD89tsZEiytu82Aic0WLUSjyIeLJCt1aW3eaIj1G33n62t2JPASCvSMl0lxYS
XKx10S5AuVt//1JX93MP66HttcH0wFhF4gA6EcadQKE0H1SmMu0CqYoKnxFqNGOlH1DqSIJcVkAW
L5wyRVwAtvbpTfJ2Pe/r5Ipmf+cZgTqPB8OcxoQjsDUZ5+BBBLvLdTMeoknjuI05r03Egzfzyz2a
/lf0ziKT1+fArpZ/51F/k34ErLTzFjRndWVzSZoqL/4KITt/9VIDnsmY0z2w3WqDreJZPP2w92Ka
u9xDkXD4LacW+qE/654USItBztIAdRRKzT9xUzbhA0pflkJkHh/Dga3q1GHSsEUSAQSiwe3c4dW1
q0u6VySOYMdnOOPavkT3iG+AWLOuJXWbDjotqxviZCLsda+S1/A+5JI0g0IsHVYc90epXOVf/nqR
x84ZdgPLB7ndRqIIsb9IBqo+tO63hzU6k10+3YbL+7nsskofZVBJY11JLiRDgnRrLcD8PUcLv9OR
0OEgUrgUhhEmEFoR15bAvtMHl4p37MuShLvCw4Zs3KJKYNPltZMSw1P4s16FL25GpRHTY54fyCZs
9nrcb+0szzRuJeWKtmuZ0zP9pnbWuV/pETjbwfnPQFOfnI8/tTuGwjCdbsKgo0Se4H0TjfibcsFj
UXdGOJUZp1wcV1Pv9B6s1jMXwbheGMNx4TZNU5vf/7MGPnDH2GqqXC5xo4ZCq+PfWZ35zGpceOGs
ZlR8/bauNTe0TNJqdurgyOX1kFLnoT1skqjqiBYvQPvHG7Lrz5Pay1YiKkBFxqt9Wh88hdnMHPwm
fxCJ5X9ray24OefhzjUvzMqDFPLCK3cPfOG/PfsFpV1V2QZc7/huiHI4t1aq44F+faOKVjWivEi5
ACyAgZ2s2Kl2aqPF2ufN9MQVtN/XYz3+2ejrR/IetSbYWxWo/TbX1KFsOe1fCkiUqI9D3bTZzVDA
0dXuYWDZ06OUP0MRw7+T4rYjgfcXcjZFpOyYqZCWxZ828/KQ9MmkKVrDIyEhR7htmqwo+ICZgOKL
mjsDHJaXfOc2bM8tAW2fGTFk9uGwcxudaV+lzfPT7h0TUSdJD1HOOHd9wwc9Oax6auAKBHk9e2mt
N3iBoRrOy45v/J1Jdj45US6vGAb5wWpIR5lw6MKIOm4QkPf7OrV93hTiQ6S+m2nRkEcbYon5GPbB
fwRoUHYG+KI/xDtB/PIMTidnsdI1x81WgMY9If49ixfZOJn8w5ZtfLj/sgoz13qg+sFxVw04trdm
3ljRy77DInhWe5HZaPVTEPqC0LhJTenhBA1zzpbcHgly98tJHpq47cW5iC4tWj7dUrKRabL/hTst
AWhQ9pO6UvjNm9DMHPiuN0NzshHvIFB7G6zo+BPf5R+D5OezcsT960LG5nzAY5jXSCV4dCq6olWd
v5hxPipTMegISLufgsknHz1KQ1Q6ul53xEjIgz/eIwMDeYHQItvbOuQtEBS+xRrgRn1ITWiwymqG
YVZHbtcjke6UygwwHGes+dNLRAKSkktgghAYGoy32KMmYHrIYii15Z90gQe8MxPklco0B0wjMf13
6Rq1Ui3r7anUe+V93/6o596RACWA+6XE0s9mS25JZaXBrOVqUJjjnb0iScDm4/VTqwtnU7kA0UMZ
DYjIPivcN0oVXd1yxJ5CzIyMgiN0sUNqWj6tGI2D71VkKPkt1SqxOunWefEJaEeynFKmDOslSb0H
p1rooUtLXRaveCzBvTG7MZM9G/oxfTGwT3dFHbStSF/wugcWwZB9CoaTS4JfTtLIDKlLZ0RJ8IAT
Q/O75eat051Nq9YgTgOHC01JB7Mg6HVJ4OxR/NdTF7DAcvLJbCFBKAGPSQ9/MXJhxvHiMkClgJeS
Sbeq4PlyBlfI/9za4icoziLXH78S7TNb2g4VTEjZRmC50e/0qb8gB80FJHmkcf/W+NVVHiq9FGOI
/ZoO90cyE3f3v4Ikjbk1EJrNilb3C5trUHjqlf244Ql5N5P/jKA4G983WxOQCWxbx1xeCrlpkjjV
xjxH00hxMoWWjVBU8yufXNXzCcm5Pqy9bVZg3qeqreLHjbH23JiZZfel4OSTquhCEoLtvPGIjQkg
gwvKPsOY3AW6ACsGetADhc7+4o/AuMbLSkCxT2UfGOSCQZ7CfT4348LFxS9hZDJqcKe0jVfM/FRN
QQNliroY0r+Vm3ckrCKsyEQpGwdOxFCWaPd80cOMRv/5waZ6tjiEDI3BjBCsI+jjS0i7K6lnJkJG
cHkueeShw7F9VBvg8oVnGh6EV5cK9rBx8F8W/DLKs/T15e2RA0omYz5DWT9/NYVw888jYZJ9GxTq
KNB5nyCoYTye8iA3vO8aTO/s3rVmMKOr33vr7gDAx66dD7UAulypWDATiHW6wsjHzPVWbCxaBTnw
NYi7rLJ70/9CX2WVCzsufm7sSnlHl++HUF/jres6m5/NL1ZJlDizk5TXINYze3BtDBqVEImql8Nj
t6h7RgZ7rim+yfRtXHt8Y7zotApsadTvGC2mkmgfxSDODS/S0Ck207BHzWDOVW3Wog2K7LkRM8yX
u6/pUtV7bEJ8Sjzw7TukheXGXiIPjPZ9BGrtiD4WpWQM1c71HdeDPrao0D2tm9u84VvTQ9hfKmQd
TksPnOsOKw+9LyHU4ZQxWjvIcI1G74DCwD1hPbiASTYs2ClUsndCx7K/YF9nHCNz1fWdNeAtkO5a
vPhafXY0hexHxRL7Qczrt4vwLJU7ufazorp7QX9AG0WLteql5PpvFcjSqGyaxjgTdg5Fth9bf4ey
1TtOXGjjPXiavymouFj+1muFQcUTshdXACYfYgqSDwU18F6k+FuDrAsTcsIm6bEax3eXCnGy6DMT
U79UoVyMSStSsR5MTYiGW67bWgo9BeUj9oOJ7ntHt8+zEcAQx8r//UQMx129VVYhK1v3vvufU6pg
PvK/5U7gCSrrwVo9OoqByPnILkv5XSGepW3lNYxG7zlUDJCveASuA24RuacSPPBOnUCABkMU+1bt
4kvOdhwfeojatjH1ZaTVWnkb13qxCHHsorGhd22E+eFrjPXdc0b7/hCvNta8MxdFrYjW+7lk/Vjw
xd8NkTb1aDf+tLtbvz7U4vmA5ufvSZe9/hqW42CLZJ7rKFp+cB1K9Sq53t53tSpz1jbqdE+69JRp
qS7yK0VXWKjJAeCrqp9iSthln96b4wkZ1CWtqqPkroWGv8nlE/WXj5x142LW6Gt6QgTLd5OC/lc+
CGTpXakZNxu0WeaYWQZVvl6DrQGCmoA1fsmBNtG31lRAxp4tSGIKcK6ZNmQZPXL10EssgaFEx4CO
XHQKJ6tBtVEu05XO3E8ey0woXCJnvhGsmxRQn7+QvX6LRbedKxjawaOm/o3Vy6xAJwhc6xbzu7E5
C2rJMDo/XNGw+XX/uF0IxmenihGOX1+oy6xvRK+CoHj1ZD5kgKgHU/cxOmluyQerSUtaBO4MulOE
+s3yedS3q7FxbYwDq7wzKFIpZzx1fQ+QaQTSd+NibD5FsnDL+KA6RZJ5pXKCiwa5oyWmJFpkUw2w
b+23KfxPghGE/a/t0UY9RGi/MCOOtS3953hvlEjmVpcKmyrAnGicCqspCExMgjRjdSQ4ZM6pYNrL
fe9IaPNryulFLVrZv+Q/Tny2+60sHZL1FQ4WzrqUdcd5jZX8yLi9U79EaGAheYg83FM20lTmB3So
I9uqK7qGwKHnybzgIctkDZTXczXQjG07TN7WUdfiZ5WCU2Jz6hxcUqtuQRr3EiVo/nO9VWz3Gm4B
5ya6/X68HXIb4lvHWY38t6eWb5gIwC3ifLQd7ESI8cNbCyuDX089jmvYU+7l4wk3ha0/dlKTUZvK
YYk0BCTqRIekH9Sw+QWPIIR3yQm5GRfFutFXJpu0vQ8a1/XyIJHLIsD/70DgU2ovqD7jkzMoVVcC
W0zekP58OawgHGnjBgEwTr9sWKXoMHylancGAtESaR7QL2np5Z/KZOO8MfIG+o6B/KJLbXFqhrJK
57T6cvIGFF+oak1QlUxVzexrgiMstydJQaOSNE3V3c03w7WFHZ9n055yKLIrfTwZZ6URI9RBa+nh
rcBBcluxCizwX9w8b4Kd1eHATaxV/kUfKFKDUcAGufnaCYMIV47o+ZvrvOaIbQl71SRvmfa4As/t
llkg6AADCqasJmLOxDFLtV/EbdzmoVy4CQ1eEagLjVe39oFhh0Xnf86alWxM2HlS2yIFRrkOtHBC
CRr1DT9lswwFT740ubdZ09SBNGTm3je/gQ7CxryZoaumcJ7KYkNvYRMbnvOCTuIS0bJRsFiBn5b7
k2T/SMVDSXScpzSa3cWkCQeZ+CtKZdOn+sQt1wf2k7VB6M2BDUYOEclJksBpnnLAyxR3KFMH3s9v
VDEeZmUR91EJOXb+WtgiGrypMHRgg0BGmUc8ailZs1v7HcN5tQ9U6n6Fg121Hkpj4IOM1CwOjwvI
+yMTVLN3F8fe6evuDZ63XJLYFLpiQJtohmk8RcdRc0shzbNag9a+HBdupX3RxKT9xKU64BdRBSoK
2HSeqA14gInWE/7Vkjcq/Oui3z7ZNgqmn7fxdFyJpQY/A0329Vzc9xauCgRobE+KiSU4Wmq+QDCp
tBczQeKvECeI/8lhP5nBRnMqeqxCSOyuwchXqHIWIBkeo+tcxqJVMOZJtgvYT69wAfD1gBGQxqpX
ZISUWP7/cURPHf/At/Wst4csVreAJtA5jnHZ8mKYk0SXJFwFmKlj2k91bCUVtlAgS09FLY+5MjX5
iXx33z9BYchd1NPf4ecbuuqM8LFt3XzPLSu21EWPtrNRl+JpZfjjKHoDuJ0S1gYiv+w2kI7NAk8E
YMo9IDbBJe3N3NiJOy2gEXZWaJBFE7jFDNfH3WXbsnw7OCozB6R0k7tUtY06VcfpaSTljzArN7hc
Kfrol2Lhf+XMsk7g9gKwqroqacveFLYwatzUznowsJs5iPoti3FVm1uEk5ePGB/4tpVGYSBQGgam
l4c/HegPI4BYRk+wGEnA5DTXj9ZIg0YipigE06r+XV5zQ6sSg1oERZ8XrBeexbGprLd2eTPaJ8fJ
aK1PzfvzKr26g6XbHXVmoWfmsvNUfvNqThESBblDyPKgEJHYbVEYNdGgti1lzy3HuSu2Po3UQz9m
CLBiqO2tKMuCuzrJZ3svI/G8MCrakGTmtXu239BC48PLr165uhjef+Q0Zony7+uLiX36j7BvlzW2
WoBSqRh/VJgIUKdf1DrAeZNby/3xdPsTpic4rRICeRvphOluxd0Pp4m6kYdHaOpT6tzG811qg6/U
CvWxHXxvcrfBP4XjWPhzZv3ZeHs8Z1chfagfLNPiO5rgHgqhFykzq9aFTfSOpifb5nSc9b4ovQ71
6ykyNWYZg7aVsIpe/KcXCfDy0Q6SXyvdsm/VHd2kMMCdrkhDdtzMa0gIjx3/QA3uAzAWnhQ3zODU
xvdOupJZ08wBUXb7e+iaKiQuzDMuX7lO7Pc50F7Ks8V/t4fwdIkPcY9NWwRXJC5ftb6sha4BGWYL
S1q0j1jyUATT+z4AkFXRnA+ZRhSU5WAAvNADDDFZOsIIUJMFtXs9xTpOqvXB9QNOmtZQAp9YknmR
OV6Uyl2OeFN6PMluaz6BY5fpx/9fTlf/N1LNU2OwXs1msVxorD9q1AStCx1AcimaMPhK0VVe7AXc
vnuz9STeAKIYsnNFGTnVOdcV3vhG1IBMYoYKRzS8BhCjovqEdU9N7/2yQrul1B/zxW0DqOqgKOJH
Z0l//kbe8eP35D9tEF9XxO+tFZneaRxINpKiEdMKYcfX7Z4fNhj24ajpc6oCPBczLGH6pArezVt/
Qkvv2LFbd6aO8uIk/DFtX5fwYdaSPXmpuXn9w10Cmmzy4SatwFdjApSJcd8anX5a20mMfiyNhhS0
JAwB84bjA8gRgZEedvBq38wc+a1mm1nGQW7Yh8nalBcCohTTCX23PZyE7QIixMIKllL8IsazELo8
/n8T5LqKsyGOOEPokQquArilixvy+U6Geb85BIl0/d+3aTMdVNs6YE6+KDLQRE5khXIXdFW1B547
tq38g0FkpmpvK8XJ7uv1ErXShwVHN6S50t+Ox7ZWrTrgDwOrOoMnOqBEb9ZoBL+fOJ1z9jov71pv
6o5CfpVTvhmQR1ThRbtf8vng1t/ZVxbIa1v0L8l8Tux/OAdiqJ1mQu4TBROkxlkPZ0S1KfYd1VsL
kxVOX8ae4IkKvHD6zSG3JrbUBYLL2ft75cJWCfBMwoBBubQ0MJwSlbz9jHXIey0lB0aDxRHlKgOK
1hSG+K6A7S/GfIVfle2m4nzE9ohNpPXJc0ZkqBnUaXEsDmKz+sb2SGds1A1Izdklm7nGTH7Wu8m9
NGaBM3fZoZv2lKQ8ix7Te+JHvtqbZh3BrbtFr5Fxos8JGm3VVvBgQbUGM0jSf3iX6C5yvir+/1Ys
rRR5wbEGC11ODqwW0FEFXz82LCKFAxYAYkXJaknf7b2tQsQDsIHnER9FiItZ5YED8/Vkw6Gpil17
Byb5L5cI1zPUiLsYDuIpvCRIteUhrNh0QCJHwo1kveyz8j16ehT92Vq/fakHxiRQcDGSVBtzAQVh
zOPWTJaAe/Ifr67X1WAxvI8wr2f/Dwnp1HzWbo4+9XGjpNwObv/3++51FBerQ09ksEBoILbtzfK+
BMmA6DuuepqqCBr18BOjxzK06hrnM3JKP9K++GWUySTXkwWCQ57XfrZKB17aO/VkzbOZAlzDOxLP
+oGfXUIx/Ekp9/wCwkaIiO4qtkSkX9K9/35YI2o+xlTizCufeiEPRMbxfhKgcwHa3DrS+d7HJ42g
M0M9G3OMQftElGKY+VbGkXVV96Vd4rNEpzIS0lP+uy68R7/yc56jG3sQrPkDBWem394seGln1SQA
ZMu8H5MwE2qu27253HUfqhZUJpPlz56P4BaNhrWecgBXSpxIZV5M47oynv93+9+dTRYHN0yjEH91
tf3ZZ2fYh7CpzWyXr8qyP24kgQrzP43nhUd8Ix7HxZnzRGB1D1+Oi1gGQ+6jjOFZsMmpwCyOcCrB
T6l2qWIlDflSP9enhjJ2ucmhyjECkKUV32pnbISW82Fb+kkEXzmSc/hD+xXZx7K2JccLVmXjXt7V
a4tghx9fI8AJ2A7NoAopZEtSCbv/N/J1aNN5yQAejwQ3cm3dHU3XNSH0IjwJnfUyo+mYzEyUrYUW
T4cBlUNQKEUUYrpUdwvMuUVlzWIKbjHJ+FIrNr16Uc8u/AxAmnw00RKXYEGZ/VMlY7Rh2Zss1Jjq
K26QavVa+IolsRURHvhiY9NLScIzVMEnZKqzfL5pujJRvH2ayzY5xEJUP9zF2ARsVr3kwRFvdA9c
Y5RNjsMNBiwCadaZDbVr7v7LeLD25R2Fg9QdlQFx3tdiKP7DqHl+7e73+iELZdn/FEoB8R/mmnFp
V6oWqAep4EdwS7PwxMnyHVMzzoobB6iXuUwwYsyH80fDvVXaxuAwADvlCEuOtI7nw/AiqyhQeMIG
Kp3Y6HWyF586PNCfV6mjTiZkUT8fbIBzaex38hQhFLqsok/09v6iSFKjLlsf8HiIv7s2qzS9zZ3R
tgygj4IcV5lGZbuJ9XUZpkw0LgDaOZDTzjKwpvzYPTjL/da6RgiPNezUxHOc2zJ3rFVkTKk1PYg9
13DAqmSbc13Lb7nVobOOlaVaFVumlG6mGqIrq7QeUHo3cwGeRGThJnFpnfCCQQkO1l2hlEOsw/hu
foJTYjYhsHYYMs1xtM4hQ++TolrZRzNlUrX+eJdnzoPy3ZE9IQL9VQ7YVFCqcMR2f3CMnpbA0GSa
5ikQebQ98izsyhFvNEC80uR4ys30CWlNXwLG8708MgdB55inUM3MWbuGXchiXv2FTaEe36rcCLEL
fUP2uzMRjfwuxxe1vGfz2lhmenPp74oevggjncGPTjoi+RGXoSwV1jjoZoGERgkFCzO7I78UA696
lCtaGAQPywedL7KFyhgioRaIOxuQvdSi6JKT4FuCXP4GcDEVTWg4TxM8l3dG4qvyNjrqnQwRoK4s
8KxLeKgJyOu6L2lcgqCaAEsQt8v28WmOWd51ZwhvzUQFD8mUkCmPABrUMj8ok+FdkQEjwhVtr6Ee
d8RFfnzy0i6L5bza/W1o0XD6ITqhDskWCUDsT93N/1asBnSOhOSv4cF+YF03tLON1DoXHGO/Umhz
xhmS6KrgPVF7nAeZbiWfkwObik90SN7S3wKC4MT0lhKZT4b0C1LODU5ZU24hXTjG4YttG2xIShHR
aQJaxcFpAlThxglRdADEojpQYl3PKs3/OhXq0SeCSlQtzwSAv2wEzgv6dTxCnK546uaxuzr80eZ/
uxxniLVp8HJJk9NovuB+CwhfHODvk/1hlI/cCXsg4E00VBML4bEScow5eGKwUxg2zqU++JPfZ15I
ho0yg0joJSSV5Is3uPIdzigUr01nJXxdgXACbcCEhBM4v+G90opKxRELDgwZsXM+jxLH0+Lbmqqr
ipShE6Inn1gACSCOnjCdCw6RoFj4a0XSEb+AN9ASSwOb8EckZd2TjgKWYCEgY+HrDdZEjIQJRIy3
i9/Icp0eYITnmB/5d2Udx/wW2mvoLZGVlaaqxhxtwq3cz43OHm6pn40hho79WEm1pMIaxv9FDULX
VgCREG7c9MA7BI2PG4LjdPaDdUXEfoADh24/NIGAsZqLWNv95/ikA0sE3/ChRuSW9NVJrSe4rkcb
50h7azVo+65aqXCDTMGwQXXFCXU9XaVDhg3mgFlNxCzKnhjAhECnb2g3oyAMEMSRNLqxas1ujZow
Dve3nx6fZ6vGTw1g1IbCSr6IEZIfxpUfmA7wNZSR9wmleR70HlSLBCffAMvtTuRKLygSHUpVnQub
A8qUbEDe6Ih7QDn9cflZGgXn8AjuLanuZxyFA74bXmy43VraEIrIKg+qCio2j3zXV88jnDOBLRse
nHtVqNHMEG8tu8rnAFmIYeemukIuejHPxZjy00ezJ5ONixr+/KSv/N98G23ocmn5N8HDRucHLoMe
Cu2CCr72e7ZAY8+kFtTRjvNubPcB50lxMvbJQthrcyEyEh7xjaaQFIw5ccozB8J0wVn2rlxuIv8q
0PLEDVCZ3OtgletNUtVssPsX23QjtgDx7gU6RqcKEkfGCZOpqhsV8gpW4v7otsRDzFKlOSqdfmPT
9CTcAmEYYDxkVkBPRc6YG8+K28e0mdpGzaGQXIiXCeta1hgygMulJS+MnjtGIieUXwiA3Xhx6OPk
uErEIQ252uYpupZ12FQHS7OqXqMfvsHDN9tgES8BnVoeirv+w5tWTZvaBOz7KY05mBaseplmjQNg
0K6X6gX5sFmmMJJ/Ygn9bjAjPwFaawsJJS7NnVqlYiNgNUQoAvQ0ZsSQnrnNmrUncjSFbvnfTTTU
rFngHl/QnI0j9tbBnBzkSFS9ALfT/5ndSWrgnYzNlh4DAUX/eWV1zdY3Roc4ORbAo4F2cSF8r9Gc
4WVD81a7xfLwNBOj0q3lzpQNhZ0phiYn1V0BNm0YCsds1xE2u6oX+D8TgeL8Q9ppOKmjTGnwosoF
MHYP5vs1c/Drsr+M2gptfd3Vmudey1Jp6A+zAfh649NNNzBJgEC4va72EMP37fAfRg84PGXE1FWA
/hxncaYPCRdccPQglFWf5O/31YlRXjYEQ8T8gEJRYa7O4y0Tr/5NzyVgmpCR9TUchg8kPIyxrBv/
CPe6o1WkCXm9Je4U06hgx+yaEsYTyOE47DH5bDgM7mzuR97GQYxij78d7+/WT0ecmK8ipPGBGISh
IawMabnSepYxp71Rz5bZbzOQ/2kWF6PgnQfChtYEHSdSvftrNsAQxp/WgtFRpUgcwV93klURyb6z
3x0rLkcZOdP7xbOicOsZFmmFPcBJ4zCCIiSN+ghZffNk4j/cJs3VVdsBFkeWJ+TaogadM7ljL0ls
w3+N0JmgjlRAvtXqvR86eb/b5mWc8yKC1eN3eOF59btQcqkm+1HhsWoi7lN2TvJYQNXRUQ1lMW83
7o6juD3gbhDMreiZZfACsgzsKVqcsc5xYIgG0L00W2ocKjnASsy2Y5s5bfV5NCjbWnZIpBqDHDYg
5n2CfxBro8LeiMF9UvXx7LTFUETC8maj1JS4Ajx/7X69LCw7gIpr3tofn4MTqLPHB82NOIgiwq92
FwtzItr2timoG+zpbfM/dtgDlKdurae/vUrun1PQx02j3ODa0KP3TgObp6tAAZh+f/RX1st/Y0in
rCjVWEP2SPtLGgY6j0n4Svl2HSKOROEqSaPslZgAmzFWitvf5oqknE9aeLtYHWrkthgkL9EjQqKe
LM9b7fjV1g/QnJ1Pcm+v8UqSMQaBDRbb6qBmocDdjD/q5mkB9qxmlfeL/wZxXPE8ZuMLnTf+EjHx
MRZf7bcObzqhb232DoNhNcVp+aqT6kbcu3e0lgP1C9puo7XfWDes/4+zmDLZQFZF4XTR4FUSAh/O
uGpUT73+kPuRGtjT3vwsCwr4g3SDPV0P8k81rbyZ4WiKQCH2adFI/p406Xcbx/KnG3BffdwLLF4J
stWYydZaY6fq6+G+2MP7KCRp89rZ/aEz1PXpEDK0JhoqH6Z/l3nnuW6PPsH66ySsgNPnsV0Gufj9
v2r1Po98NJHDV9ol36v9XQZaCprHWbTrhvEy20pYbaq6Wp6S68+8yrMJa4Q00LPXJuEkPRwkr5ib
tXzrkVgguISgCIjNvP7gzEDEpBxgUDtr6D9K9UJQcR99yk9CJGAv2Zyg5T854czPVjh1iqF9QbTB
oF7+f6Sorr36VRju9iMSDVtEaasCTEn6oPSxviwq/C2jEPeGS6pSD165pX/ZOxq93E9SRTJFdj9k
2kWTGN6y647whWCJv2L8yspgoFW0rsmxfy7kyFrMfIRLGejnwW54ozywz9+F+Ztv7HlaP9IZXqFQ
9ltCk/16/Gtv+GsqUW4kwyRkdqDWrMaRpBN/WM7DZBRP3tRUqOufav3ap+QubHEYcDvCZy6fJf/y
zcXPcXiOqp/K6n3q3TQYkdQbUUsvXNWWWdilIBhHnC1hJIGHOtwGMnwAXbep7DjVtFQsf/jb7l4s
pUkr/KjKQYa/3mAuCu0SHDKO8+HC1Tph1J6OdaF4i5E6ajt6Jha95veS8Ax94zo0wnFMkWD7ut3U
BbLlhL8tALsjiRAo0OWi3bvZJtNGkGsvFCzb9i1h/Sp+TsL2YZ4RV5uMFqSAnZN+bIkx6ODalZhz
GB2pStJgpKh1zlyVI8FqNtdZ0EImeJ2NHtxK5n0C5OdaxuAikE9XL3MzTXuG1T8qy3ZKOm9XNIKr
rhfXCbVLuJzMhBLrWgaWsopKpJxTUgKmW6zv6jb1mJvPsW3Kmg77wOuoCbi5rlY51qa6zlOjD4Ds
y5LRQeTDsNGxnrOE9A07FwXhiMfVEdobpFyPUQ8z44a2qVSZlnwUrtWfLrb8akQB87l0zVCrjg1k
o8F9Z3urQ0c3HGiJy5xphbvjG6jrNpg9U4KwEBeemw5VIOra0InkQD+b3MR4LmiQd4GDzsEXNHLH
vcLu+0mF2+b0+3VxWpBk5TG4slgDsfjFdmzcHIUEa4QAzyKvL4Tye1vdBbRQ6JDWi3r+ceXVQj5X
FkRkAH8cs3rj7myOA0qau4SNesuPZbhwsyba6kGnqI0tnKmXdiDVv3VgsTwayJqIAC5kZluOd/CX
hEv5gHTsSGmhQ+Nd9CnQXOH8OEiHycjpMu83THNV1s4xmuNi1mPdp0++9nx5qY6oevuHLdy8P/el
312keRkhvl2FjpKNZAUIfZVzl+rX8y25M+gQXmuBZwl4NXJCiZSHZyNT7mxI06AlDBLVWd9zWkX7
7RoRkVpHqfDjrit/3W47RyuArzr8KWBASzf90sseBxEcmxwpGcUqc+3IRZFAARnouARzXdQqWxZ7
ksls5l4keK1eSdvYei4CFgQylO1sydkYW0vT+TX5G8bJ4M2GwYWKPLdf5YYdUBBJlnqYcWwXP7wc
j693RJCDhQol5tfCbyveA6xi2BPT7/2+3oFMK3zsJAWOflSjEDhmsAe7jS7SPhD6La9lCK7oY0Zd
aAb7mCFf9iHSHR7XfwOjjzhxlcR9i8sO0REc7giH+nwRpQ6YCPgW/tnlvPMvPgy20V5JiUx65bV7
wbFKWD7fRKurgjQ52gHqSwIIw0XvDK1GIS/iSTC7YRvjh7/1U7GMkIgY4YsIXhnjW8LeGW8BHmNM
sDliFCrAFTIeZj4pHiydB0QiQ9IHsRpwsWAnNcwPevNAhG/1Ru3rly52hD5+19KlT5hxILP6Do+Y
PEYjDSk0l66ZWTi00IpEYVYoNvMwMJIdNuA+AUJSFS0ARONIK9vaxXTbFZYpujYf0sprIDQQyK8+
OZgGFBItQBLqI+qhLy7Gvggx1WxHO6JSjG0LNYUMFzAIePFlnkxNUVaRt7HA5oOE6BtF4m0sHn7H
jnYNMcVfo+w2Ryn+mml9KJY4c8NhW3x8mfBDbrJChLbhxCC6g6NbgH9BsMMA0v7VvAOeMAdSV5zg
UsqriUoq27B8MTqtul/SXMdfPteQr3hZk70F5frg1a1GF+2w9tGhS7ztgMZShpoSDGjgOihXtsMD
x/h3WVxmeOpTkioCKm21tPTZvzVQqv2eTeCBtaSF0GvpfVbEB2/5zu66d7R9beFHX+Bdasn3v08g
Dvu1ce0Nv2B6Q4d1calZ9G3fFcbFeuoPLNp/HdkcZMuQHAmRjKQE8sNLrpouLTuNQJCaSVlWlVyz
71kX3YlNJs04I2MxgmW+4uBI9xOSzR29fOKZFqy6RMeMx7MBFzrFzYY7Ze68qitdluM71iXIDs53
DC919l3HNAjRIsWrX7tarEGzcldDOHbcT44H7PRAzfDhlICsvK7ZyOS/TGOVIjBf635zPfkHxoul
YNoGehZVOV/2Q1rctdTF0PI7SgqrPuUjcPvbU5mm7PYwXDurfn9xli0IHRaP9REYrfy9eJIVQhtq
H6nhLmQBLSw/0ppdw2gUiqTo76Fd19REmLokL7xo5wQi2n5JwAkz5HbE13ua9PWdTXr6A5bTNWu5
78c5XbrB1WecsElz2L8YJ8uN2bupNtlRZ1L1QzopsJ5h/k1n7W+Jw2Ew36SI4DB/FtoJzqtG9Nc0
GvU7LpUfPIkWCQZFDEWbI/8+opUxTk0obYZifzxA2veoNHJNT+F/EjbviwMVAy4yDUeUQ97SFcU6
3EG896Fi2Tn7clrb+0KFbNh6vag/wJuPbuMS3hVZWYoxg6LlrlfG6IhvJJuDiRugRj/pkypskIJw
eW6YbF9/H1LDyCEQ0OhLtT57QFCCc2t2yVI62wQISjiN30PcK2FBbMVTSvblymyvy9qQTF+Co76u
/XZgpeFgAAJAzX/q6AJ03f4q+DUdb1Cq/40J2xAd3tsKpMADEdCNQ0z3/mh/7Hdi0LcV7KBrSLe3
cLM99SKRZmM1a00qMqXZ0LHJW+MOnR4pzQMJvnRH08rUQHsiMm+nB0tG0eklTj9SLIbWyBokRAfm
CnrDo/L/JBEHnZrfjfVUuAC/4MlM4cwPUxI5Xp5spzAgTU4Q88FfDyzqGhOJKTvhG6B79+gg7PdG
vqwEY7Oc3ReE0vsDbFxjvpHq518zmnKCN7+r62t+HWezLL60S2KjBubavFLSorVhxf3Hh02oollu
i028oWhfoPv+MSM11KuBMEgF9MSj+zGnA5Do4fm3x+nFdbjinWw9swcTiQGAgCud+zl1YvyZmBXE
dwziU5PhuGllidqYnoQl84dlSMVfCtGBfNyl0lXUpd8DVh+2qThqAC29/QHtctfdJZY7s1q5nL4e
e9Ujd4IipeZNSM+bATEdiUSJv+pR5MdgLqTTK33xA2Z1e1CTnravFisZXCJCwJL5+qI4cURPUkP1
zkSHDAYUWoZXgqh8jjr52ERL8yhMB9aHpFAcU/zcEh2zQmYSfNgsugrUghgVBrq4tWAvpAfZtbDf
mY0bJd7oq6D6kz8NARfdVt01sLynL3uZGlN5Vi8NC7j0suu6hODQtCIjweHwOMhx+URQEivHPYRm
ap1s8QaxcOn/PWq3oU97wYChknvS8V/Bb1KJpwittViZitdWDCnNLDcXSafL41a+PmYu0quqTSBK
tHvv4I/jD6L+16Ll/eYAc62IKttW8jIDacSicTmd0jCS9HVxRwQbguRNztISPADELB2xs4IIHUjQ
fTW+6UddjGC50ptdKgN4SQ4mb/9OpDZCIi9v8A9eNOs8DCXbfENYBTHrX6bl7y+Asgvi/17kiPnB
WWBdEoXKrJZgqjLkbiuIpXhIrgdELFcTHWx/QuutI127qg86kGf9DQFoWPMivGAVg00kmhqA/+Vt
nW+5DYr8pwlQM83YCw6dRAdqnr5NeXyF9cOiKnasy6PdAS8yUfb3PSXc4PJXNaNTC0qCdtH3R45x
Ltm55mRol71PRmhBqGM8C0/fNBHlWUXPW9lcJprbGDC9TQ1ZKQb0+uV1kk/uljkcdVtzFy+OoO9D
v209C17y6R4gaNohKji4a75He2RRKvGtiqJ7/brtmhNM2E+6AFKowsDuSSsWtoqjIacpK8cOLyt9
98QF9BsvUsIPnEExGJh9Tau+SIaSIcDgCGXrjUQBuOP1FK9rBhJzFybRcWwWDJf84a6Gt9JheGUZ
koTx1Ix7LSdACL1HWJwhRpUyFryodpQQXWTBfngTRuS7KQs5eeU635LwkGFnL//Crtgl99M1z+5r
y0aFKGWIa1hysgZdtBBVEO3mXDa/Ws9a9kzAWIVQkMqqZXzEPL6UNNc/zkOFlHJbt6vF85Ub8W4R
e7ZYPx3qNGUXNSoK9DAa4jAFFIQBaDRDPg7+9mH7XV0RsDivfRRKcGQJoGxkrp2RRZ8X/quSkNK5
XSVC7r3bg/vP2AphFqB0KRqM83PRmDk23Xvs7R6ks2sEZyzPsgZVCfISzrRUISbzOjfrn3gBufRw
BC+NbWHW/0xG22v0Bpfu8vX9b21W06G/BHA4eco7iSVAm+jnZc17OLXash+wEJqLRS8jtCGlFmob
k3wPGzfn6NRdu9kSBSj16EjAZ3vrcF/fGV2Bf9CbFqOrIKwoLx5fo8DNpJlsQrb78p8tdka4yd/v
WgcQ3gdQ/L3USZLoZv6rTY/jr+yzfN+q9TRVo1K1tARx3M+tBaIJT7oxwCkIjjq0wj1Jzch0LhUI
wqH0oII74TCirWs1L9mcKNXNeyy004t9EOw0gkWRX1lDugVcuDkArFJ6WfYlqIUI3FGW6WFJK41b
ufw9Z8tvBwj1nwShjzWydLy8jN6I3L1zks9y7+6Cy/uaWDZNjoC0CzHV4enbtzhmJG8NrP1lUUvQ
ZtNYGXHSKoro5AiSWGgJZSYaegwEpzeSIIm+/LfzUSvxaeTsUF1psRJX36nDuyAw9ZyeH5d1Kyqo
uaYVhF/E4DP9RaOtJoFcumuLoyzWf0AQbvBulJKtFTmDmZ2ddQBf5OOOUJ4R5szI5QooKGDXoLyq
BkUORoCZp664lgq3BVssWF9l/GcTmbJiI+Ku+xODxCiYtLTf/tPZB7OrPZStdvIkXCe+QvyCAR8B
5ImLG4AUXOkTQSm0oTX33Lb491Awuu75Ohtlvob5q765N9hfGijcddSXPrceVwJ4pdzRd3P+5BmA
eq67L9hz8OysdwuUDbQI+h5gN25IPoy0CBpdDzKQklDKkLJc/iP+zHzDjzvJ8ATyAwjkahCkfol7
Soq3itxOpY1ofYzpDpBZeZ19dHA8YllN2agbbSr+y6wXaLnb49JnNQY+kxeg8GthxuuVKnC0g/DV
nuqlflGOxRm0bv/CYGbDsJkOwzKIslBzNPN93M3QVApKcybxNDFmWK8d4T3rPYgscw7brxHaxoUQ
woTKRHAI4xZC0GZO2s+K2SeWva2PkKCVxIW577DkhYDCkkNisvVhhK1lTf59M3wazNF160k2PJyk
K1dEzW9Vd89P61H0uHCKBALqfHyNcwyyZhBFlF8VtY4oGGaEtXe5aSZqrOCzrqGHO/wN52/Ki2x2
HgLAT5Zfkjgb5HjsDyQEnG8d5Jb62EuVBPOw+bBV7Ruupkxzros3aaZnRUUgnGYJTrNA0WaJG43f
Po1nC+X8E+OvheF7obiodF8eM2pxMnmLNK00WqDsbm+cpvoC22x7Xe9HYif/SMKE/5NMq7ZRAvfv
4HjYHqUuCnnMMEq1FWCuWfTcDhRStBG5ujnhnRAWOm8xPVA0jvdO6R7jpDaeROaPB/NXXrkxVPS7
p/63po5Lyhoc/h9Lhxy4H2m8tmSM4RYAzoZ+6Op2gLLikixRate3GgohPgJ8Wes2V4mJ71XHBQrj
rj29xiZXSQeOwQK7MNC9mYEI1RW0s4H/pndAEWlGAyjhgiS08Qq0jBKiko9xhVpvK1h/DE+eNGkW
OkdbAun7Fdl3++dpW+NWXkXvbLZDNSEjQnsdfPy5skq9n3MOo40I1L4qWO4T+O9cez1U+oltvTDa
2Y9L8Ws8MQG7073UxfOc8Rs7V4GFK/9aLQJ4fw2T7bJ35BKOEqxzd2ki5NZt2YylVxpbjcjuEWVJ
9G7zAzgbewY6IfvbvrWSaBVMlv+ZKa5Hlj8Jn0U2LaOOr0hhg4sQPkB2bfPjHidBlPv+1KYRYXag
VmhKjPzIp/4P+FN9ta1wTgNgLGMjgTZnp05GbiZUlbnRMkmh3qIoeUDgtxdGJ1IKVtXuRNIy/U3V
1E2xC9qhj0PMlHj0P7h/77bZ04IR3py9A0/w7CNTkAnIyNupUOg935lCfwT1nnxEl4FR3Eqaa2Ct
NWtTvd219cn1cRmeM6QTTtblmlSTWD2DP8gutlKLJ4rHmS0QIqRJS/1hs5PbQ+O03cTQh9DMWjbn
Nq6QyGpZcr9NwGds0WOSaBzLahyg0CtgrS/YjBt5IvMNNYhYSXX0w5lC84uUW9WOO0qb0wJiDgcG
JbyidLSVdEXCEHfEQxxDA7s4RTgtwrsWNfaWV45UHS8f6JnM5ViZKIJ2VPuWffJMdSYpwPhz6dkh
i34wUKJN7l7nXwFOWNOGGG6xIKU0gnIWEdHmq9YTudP90HR8QmNTVv6OKlEz8wGdzdS4jHzJxE5N
gB/tEX2TMTNcpMSBhWfvpk9kJoo6ROJEZLAhB5mgYxacZTL2DKUVggTCXgwmFrO+o3NHz9vXqNat
Q1Npm4GjxO+uDgCFh+/M25CwTC3u97ArF7qnQBrbM0Sb7HpzGjHaJnTbqELvwG6d1DcujqSLjITR
2ABszjAYAlNtWYZZSrmUkNPJJZC7ODpcQgKP6jJAoWoIoiUJ0TQEiIfCvry6Fd5e7hj19jFJ+kHN
0F8WDcOPNvg2WaJCZSkW7ygjZjmzOcr1usDW2KX5p59jNqsKDZpvL7gkISqM1pXMmkLdUJ6gstmt
52PV7qnw41M5XxWwlsAdXsd8p7/D5bRa2DKqvuN1vGaCaYnBMqoA1nxwro0E0zlIf/xNCUCgj9MG
70tPqoumoqxEtdxbSd82oHCsG5iuCXQqhcYuynahVd2fRDcIUanqM3XUWXtKDY/7bt8jK7KjymyW
qpmIk+NyflmPnX3USyHONgMk8XHizF8fm1JuvmXkmppvGtAobGcTt+QVXJ7c3n49k69XGsTUrbG5
hqYW6gq6KZMk+nkp63IWaUw2cOvvKZYh3SqunkY94cn51e+gigqRi69XzEjcZBasjWrCRWxMXx/H
eU1rarFyBSt2yh89HOiduH3IYRHKNHVOzWFUJSKEoKrjxvopnoo+0N3LsNKvBiadMaJCxK3Nnc7K
2QdRcnuP8RFp8ynVvNdJ9mI2s39PMfqqvDuVTJ81oQvtXdp2Wau0XL0hekqSusaoXyITqucJsT7h
jLtjRuDvUMRHnjQBCGTYwPnExuIhJmmTTBULLa0dsPK8X6QZ6i7rpBIChPhd5QsU3H6WPn3dEMw6
2J+7jqFEg7i31F5yCAl4WilzGWsgTsczDHe1zXxXhbTMa/OiaDdjs+i2myL/vqjoFn0s41byn8PY
kfWitt869Ts9cM5dIq2Is40mO724+rS2qMqv7G18wfyAh36snA2GxTwVk+KWWCTMOIB9wdChNtkK
Z/7DJeW4b7uxzoJK0cH70XXAHkNi4dGPUsSuXUr+tdbJyV3WRmHxBUpFP85EKlfseRLrhXSnE7M3
SbS1V8KNOyp1XRuqSclo7mdyHGAbPlJqebHaPT2DZE51XRDXhJW+f3TzeHOui6/f3XAscmkuhrg5
X/y+2llq1jbRcDUTAfHl1I5iyu3gicnpcBcx3dskaDR7qyka5+P8uHbdUuZrFr3Ok+T2AgBCXFlK
4SucDDe2qztFzFZQlypXRtIQPnHOuTAzsYRcrLmf5jZMQJvvYhBXXeMcx9oGYps4Ft3dtH+2M+0w
feozjsFsFXs5t2xzP2uQoSPeerZx8j+gC20u2je7w9eUjnSH9Lk+6MFllXf5/Abwn4LP740kZDzM
y6+JnZLRWypf4v1v+sZ7fEnbB8GqSGIt2nua/T8KQugk4FbsCb+DgcssOsOZugAoNR4RPYQi+B89
qeTCOurxhmYvBWP5bmUnHwcRLfpERng/cLQh8QigT4quLUoG3Cjbh85miuz/GH3cQkOXIhWayA/D
BGp4FeR2Rh4gjvmXqe0+BrolF/1T6sXGYCW3TALVIWCe9oOraxsxKgp7z36biSkvlBY0md7Mfb2z
UojenJpEL8u/7G1DLs5tSJ1NbNhZ+BD3tHbBQ/Z+wcrXrTqaAOeDAxpWWQEZISqE7dhqvPTh3THk
tVY/otfWmLYjgymUlQElQxgGXwLJSeJ6b8SFuK2cpcwWi1mO3ei1fescrurnXr15hCs4J7xyPUyH
fhWWAkcC1KKyPkSGuupPS0yIUWG7SuQ7hJI/BqrsC0Ndgk98dzIjal2QyxDyv7IWeZu93plnw74B
2M9DO1xatT8aeqG2j9AWZfa4Lmr/qGpMLenKbo3awh5965/XCiQl7+LrsLkGjVIlsUCyMHzAwR/M
QI4uAKfjZUqNXTVwFCuAUW5YX5g9jEVfalXFVp5vd3jWGzSRX1eHnvFkwzJj4OWdt9b3yKY+8xOP
cMgMj0KfvsVe8buDQpxs4/RHj7lxVxVqsjmMf4YLDYbyOfyglAe40HJzinMftk2gCMAdSQ9JJMTk
XRSFzrbgxFYjTVLJy91VaC4eTzgIBjfKDL3aaOOpr5h3S5jRCKQ3AWQGSON7qfej2fSfuGxriZJJ
WwFL7hoLPAuvjeggLbTTJk88baQBVqJMahK81woQpAoJJNwKotWTvgYt/aM/tKboKwQZky9hsOJP
73CAC9s7q7c4D9StNdFeGG7WkX/NozL+YNfjJahKAG1tYscWppqWT8s6mk6vYkMXurCIfcCfQuC9
J+bogsgpJ+vPaatrtnAKOCruNZdh497ryz+mwQNIRUAJC18i4mX4qt+MnHaqjw2wS8HeRitUq42z
z2czct1veCHTbiWrsjXRTxJnWYOLl950/OetBqQ8qT3Ls81HXbGWFB4c9oEok0bqB/ielG1pKg3+
XPYQFokts5RluV0FTgT+GTQC0K0KRxEoqyakXuRTdRSWownyVsRab+qM7liC80p29csPO2QUwh4I
Qgw2SqR1OPtci0XZEENySuGsgvlt1ijdHX4ftHtJZtB7kNVObJ6Fo4d+C2EZ10wq2ohr7GhvAlUI
Miq2+qgHoT1X47/SgWZF15fi5JSNe8AzlsG4OMzsNRGGyFLRmenjxJDi/J/cxl4AzU1dxyvpm/XL
cQJVIBrHL1w3GPDxVzg5MbkNqgcaHtZNUyUlUtq3o6yzx2AwS6oq7YAEfjobhawAaoanxzbkgmAe
WBr3Pb/8nbmbYU3PUomWbNNcNle5STcEgfckrWANRsCPAC8Jt+fIwevtryAmJmFj3AxRVM7zzp6l
LovXsu6lolQawhBz6SdB/A0eBA4y43fX7pzq8pKW53KnM8Aa/3PluWFqysZKDJd4xC0KjT/VYjGk
H+MrT7ivVbzaey+CScfeEcOQV/3iUA70btys1XDFFBgkw9prIluquTzyHBLEp71O/7AMt4VRfuBf
4J0z9GffS66+6H1+eWAb6f11BrWYzSrvG+0wFHAmE/MG3zKi8pKI0/5IKAlZTjZ9vaUyMMmkiD7J
PADBpdmfPKbQ2H4EjZK82Go23Q5um66iXqK8AVmlNqbOBk4J/US92DcVTEmtephcUjQ6tPcuTkYd
kLSsgYU6UwNW6MANiyAH7O/MGPLjbVNBmf3HB0ITVApWGls9GpQPtBbfaFE5rHdU3RTki+MKROCS
3lYf8XRc1CxEHxD26+1Vg3wYlYk3szbWos4W5u4ZzDbQk+wB5Hgd7qFJXCzIhcbSTS8jFY+TCBmj
0qJzRbC4utpypip8KJkYgpVUYfySURjGDyVIhsPnRTbuxfdisi9UlQGJbcx2m8da4il5+/fKHugT
3nTUcx186qC1N8iMc4JrOT4JBL6V2zvYwLz2fq0+y9Oa+3sJvhSovDzXh+uhdzZMLr21osRa9LOn
ajS5tJKFB/kOSF2dWJKd0orV+9rKWdmKGMho0OiZ97GsJgneoVB70Z5FmkLw70MwmSWzrK7buUpd
7/Lz/CBhCyXZmZy97xGgcXP3qwOBJyxS9eRkHqxW2WjjOi5HpG1z/HQIwWBnaYDjaRGmqKU0yF8D
YxZoGcqfOtdtdgR781wCxTKvamxgJVPZ0NWqtTjtd0A7vdSNeG6CkXIUnVCBM7Sg8GnJv5D8V9rp
7SCLzi6qT4FyMreffkxQv2zRLJIiqr9xAD7jgq5xnnuSXq+MX9rClOkqnjYD6LlmljUA6L3NV4t3
8wG9Ww7kLRBEgoTgOz5KwXOsmNVwWB1lVWezqUXB9tovvkBm90egC5HYT+YXWzNwRLbOZIEwQMZB
vxHBMm3jlg/P0o0eCaChq+VHxl42JkTr+iBa2Rn7N+WgDeNalBCaMkuScdKk0gPg51jOi5/b0hhQ
53+TQOrmYq7RECFeaX4n2PLvsGO7Iq1lUCs81hvbKqc3ds3YegqQLyjQWsaiMpSQdtpXyK+mcDWw
2WnIOASKC1oobbaM4RgyjssLi8Q84xgyUJDOTerTLDBCoMY4nbSY4Y/5mWMUaAsYyu7di1mipzdH
Q+F+vftaenS7ozOpPritATID2s4tgs3BcnPLaHCKRi+xsfQ6GKwwHaD05d2WpbmJ3fZLneu/6+t7
AHXu3Axq0zcBpP3cnXvcCDUWuFZFycNdWwkVd2R2q0HQ5k7hn1eW1cDLMCGhJiWvy6S+UlX5R3wB
49BfAKwXcyIClUGrX1I5oslmhqSgYtbwk0A3vs3miPBLhjvgr93q57ldU4j1c/BJMbt7N/B5vYM3
W7/omh+AGdgtED/a4wgXS1P4dxVKANXtIxUrdVtJuYgkxZrJJQalFYSip8Rl0DuwJNPMjJtx/xIP
UwNjtFiKMtl6LxjA9pxAvFXYnqhqK28VWnd0oIH9iS28WuxNYxQMuq9aPe92LqstZeNbvJTBtVAD
fvJN9ljqFJVccgROm+J1e6Vp3lTN68gIJVrE2Mgs4FOTieuXztNtQxi3srJpwBZ4Y1pvzWvVGlnB
/PfPorrntDSGWuwkxFSc9/VC4slVZEBjit5/x47cS9t4QMalHCWEpw9ECPsTE+8DsHv2P9Qh7qq9
plg9NIGneDQCmX6SLtQiTsHSYrGkN8kcSdupMD+1cv88+00p9saOs4ktqNWvotwDsrrlJ40rCLbH
2KNHbOpQ5mZknnwStbOWjCdzHirBObnE9aEM39kFSxQgu4GlMK4mpBzP1MKH01l/O9QWAjbT9bZt
8s2Ep2PbFBbp4e3ZVC9aDu6hpPXFw1IWhx1YdV/WEL49zBe8E0Ubo2jSVJfySpGv1xCDpokwFslg
AYG3aRmyxpKV8eAwIaY6lpF7nbyxFuiBcigsE2mfafFfhRH9J+sZeExxWTHAC0Y4rWmmvigcAA+9
xe1OkB1eEqPEY/7R64Hh2avQfJU5GAchu5RFrjD8nQThOzuAqELYBNmEmQEWv0gLO/Dgh+cwdiT/
GpuEH3+msbbqSKanY84uQpNQhWKLcAOvBXwKWM04QHfm/PSuvTwgEWmObOUbZA/WPmuxgwgLgsXU
UU1Bb43w46ykAsGoOsHOGcWD0AHu20fhXfawcuiQCnau92ISTrG/NBBzpVhx5IEIeTsn5qaK1kNv
zj0QaJ4VUxGEVZAsCc6LinKKXVPkKcl/I2afpnjOYOnbTj1qR4nkWRilBSSTHR6ToEqXnYCBaLu9
aq+d0/wx6r9jmThQXvmJFJirCsAsY8CZzsGCtfsmwMS1gehP338gsBOP3SDSBx7v0SkFdhbmQx0V
I8CGKJ5xiS826fv5t6r/sBRyKBcy3PHf/dIa+vob1tFpJJgBV1kw8T33dp2evM4Z9SPMo9mSd4bu
DkfL9C8fzLeQZB+rvF8v0fHzh/olGgi8C1+ICx2qPRyWQ2y6mWDOKLrdFwUqVhi0OLiewIVZLLOJ
pREnixtcrpLAsUftACTRXQemcfMi6zPV9o+bhntWD9dt67Uag54dMlx61swfALo0yStaoKAYL8Hy
gM1YY0LXkH2bWtGNfc5x3YkTd2wVCnB/Ev6CxTI+j9Jv33nfgLHDs/IXHw7Z7gWcxx6EjDQ+/3eF
gTnIOHLmLa9BSApbPWsdmNnA2a7/Ww0n8Sv9wyIq8XNdcvtpyU982XdTsn8TdlDKr4G8Xv5hhTYb
5crAUqZZ119/bCrT7Uyq1A99I5nI1d8UZjw5gBAmMAcVVm6VAZMF7RkqwJ0XcjqTG4PG8gBeG1Dd
2pKOt9UsCy1Dg/M7IXKJE8fxqhHNMfO8rSyEXIdgJpHguENHlScPIi+3pspcQTMlTwrLPMIwkyLs
LnEFBYvLnLG8u/qkrgfPhyqpASKhuWV3K1Lo1InbSoDTSrUiqBgRIsYbWp/z+lJUjle4XNpzONcz
PWLlfo/1wt6bRfuUCmo3I5zXMLO6F94kfWK2nBRcVBNY+AoLniY2CSawLqiXia1h9mkfYq5qGePF
LtRZFg8rHw8CRGh8/pnfS5Ng2vFdYELPpU7yEKrHhNG055uoReCn7wkjNnu1PH0+4myh5apKCvVL
6UUBfrNm53O3Yk9mjs6SKYBtJ63kg2f8Tmsz5xuJKzNN+40xrFnv20O7FSZRHHdNmgJOjAmEgR0S
DU3Dbw5UPZIrS6UjHN98F6Jl+86QlzorHe1fKQlBS3fIrGRNVfqGEv2IW4xAARU03fuKekUHJZQv
up9v/wdaI6GTyHr86P1VgSNd1p+fErZxk5y7IstNmsSUrxHiGI5om3VIJ0fihAWIUv6m0OHzl0bG
ej3+xE0uIMBD4HiYi1VezAcxl4Q9JOXGfCZ0nL6dO8HEHlJX7SI3XKalNLIudwIyHPbq1uFppJ7r
qQihGWBa2B6KOMUx65MrHq+vTsYro/YpngmpJyDfzeKOM/mWGIJjLXc0G3NFMI8DvT261RJB03Kx
ys5UOTjqHZU3l2Fo6F0k37fVnk3NYP48ojqW4H5GrgBwkDGEWVSPZEatkX+2fDF8+PqhRofSTAUk
1FeIuNCULi2G+u1sGUV/Fi1SBXoX5pfRPYvUAWv6ZIAqeZb5JpoTQmaPDCL47LC2JKsqnbyNshWO
UviajnAFYDeT5nbEteksY+mRCGgRhxSEAxcK17luOLEiDnhm2db8RW6immEsgc9awjx2BFFXmLFB
dTT3GiLfk5jqo9M6kwdXEBacHiDhgilN3LA/wFLh/5NgNQCGVXMJixpC8dYlaUPZwE7fznzXBKrn
jrgdSkOolsDDj/6HuJBj2aBacm1uHreXO1Yv13JxthcNIE9oMIwwoV8Sy75ghxzoj8jB8XfL0N9v
voBJDkzkYvfbUOFgwru/Ge5GgJ664a0Op137+4tw2X6rEARLIFES5BG54i1jrgq8xAK9Z+shmCuU
MjUBK5IHk8DgF5nsB7V+Y7WuXTbIt4jm6dVTLxIEYsmjzz1fLD22CSQZvmwE1hT8j6KSrujQYLLf
ux+qKZU3702Uv8iZwYVpp1ZBs9F/TEXkq1HlgrAmGUpZB9hnSOodPnbX+r7BS6SkvhFIg0p7JAnm
e9fJZJ2PCDlWmyKbIRR6Sya5YjZUccK36w0qd36abG+qUDYHive19B7MXrA6PisS+yNBUPDqqKNL
RJwef5n5aBAhF7D3DHUDdz6cmlhes1q0Zoo+Bo/GGlBIv0Ir/gTf24xiZLmgYqRoJalw4O7E5BtG
Th2gxgxfF6nwi69ghmRYQbzdGMiH0+M+aX5pSbSPkNipNNR43vDcYBQDYXNg7lb4aGVi7GgcHEAo
z1aqHykmLhamHkP4Pd0gt1iRJZvvFTGNnIzrGKLCjst46Mnfm06c8T+Qq8tJOZ3cPgAHQqo5ZWKH
Z8fDlX7KF6cir8DZVkCRPq1NN61Kw8s9SD8kindOpyRTF4MvWOKbuJ58zhx9554+CBxxUXN9X6IM
qWbSOiSML4zLnBJUbuAuqrlPEOFB6uP/yk3B3n/LQUs/sYQdVzfviW7TesxVMbmVpoRwYWvDR09Z
m5s6eRsSAJRUhdQ/Bqb9N/eXgHd9livBv5d5aTJoueKtlC/Q10WTv16yQjiawVpQ6p3FUZf4FPUF
mbjb+j89jrF/Nr2d+ZkTvF5T+rxy3dbJPhnHU5VMxFxWDsvCLIu/+KtWu4v0dv0q04/1qqMIk1kc
/1zUxQIL8QL30HnvhbESLzaJ09W6Y66pJqZq6n49OWukFvnCx+fOcVeMil5WnpCkXj657+hjUFU9
QnaCObfT9fIZdBADrokkF39sFPoco97SUygWJpf+2ljN2BLqWVxKQ7Sp0T1sGGflYRyz010IPnUW
mV1k7Fm7jQkkugn3+T1JdAPW/dok2frOUVBgpq1Hle4ATJxAZnHUBZa/wVIHztBv5o7nQiz0cPsf
s/yq3sugn/gXDRsn0p/we4TkWApBmJqBa+c4tvoVZTA8yrrH+QXsQTGq7q09M0f3kRi4d01QjUJX
UvmJbTkKpXoBGjo30ttJx87x0HoIWy0HJ+pRgDcqZXJ4SQB2p/MroJi2w6+BqjsLQeaqHFjt23Tr
vSl0+uH9ooHOJT4Hzhdo1QlTcxOQjGdTxp4e2avb0j5HZLs3inS+F9+Em119tcaw6hdv0muWhsaw
kjRM8zfhS8jxyXebH6kEE+bDKaZcExnwqHYNv6Rvpalvn3RRxlFFDlK+MmYIln7xpkX/v2EfJEnx
wRxJncRnz1NGsDAw52Q+soQNJ1vYwdRpqcWhcqKbBNwXyaIgpKs0dedZ2Nl8YEHlLgHQzLpiQUBT
9qjehEvglcTm3mwvewuYZE2glzMOQbwFItBCJ0VB7XNIfQkAguSwIkappTZmGnEYSHE1xTgV10pF
K3ZheUDa34doPMJ7CcCG7UNK2paOw5tX0yNm5EP8UQiA2HqJsO0u0CDnCTZuaOrdj1CZohNWMBc6
GT7bNvaPgM93ZqxynRXNCEIDgRudh6bebigPRid4j/JMTtBL8icFlOwsfnNwcJM0iCnrjRqMD1HA
i7OciD4hMyLtN7DQII5uYmAGLa1cuYvQXYbZMwcXX06ueEtfs/AVQyYHWTdYdZ/l7+yiXvSZw/Rj
3uddx4whlGZOgYsdIuRRgY6e6Rl7wtgeAPD9i+PloC9JFnRCVTJRbhKbjvjDzIqFZrCNRrocuyty
nWghhB5Ep9NCu5lu10VJGSjSYep0J4cJObqEswoQNygHr/Fx571akN1d/tEu5hipU76FzVIhpw+B
FMKYDvhu833fkp6xqBUStHvLdXnyGUJOvb2xzIlahRmsd3OXSZ6beKhKiOXAMfb+wXMnkCoPjUhl
LkBpM1NlwGSzAXubKxViVxAt+0+6CBmB3VpuOGlmRxV+/d7TXH8BCkQwBTgOPTH1YgRQ0FxUxDvu
a2EO5qVuzcRdMuDC7QUE04Tbv0Opwy8pF92rstFpP0iI7/TChdCKKhovw6GMo6HVeKyi87vzumXa
2ksLQS9W6Yo3hzE5ttLsmbGnhx7xDNwq0Reuip9qJzheUvN9sRJlKZNswiwnmGXkvq6t690mIZnA
oBXuM9ndimbSshZkF4QnqMR6gh4ojZh/1refPlFCouF/+ok761jR9K9HlOt8kb68CC9rOX6UVsjf
KZDdn7jo8o8mvD7anhXTLe4mtWDf89gZHQuVQDa9Z17yDuxYSA2jL0apjXsGIMLdSqjqdWrN/nYU
uyIm9IpPbgy54b8SKnbl2HTGJIX7V7RcKCj/XkPIfXo2u+Vd+4AEzPthi2W7wE74mmjo4CzWITs4
Z69SQHF1d1B1Uvyhv7yGQihxa2aaA5m+mGXoRvMyxYOkEM8nf6kwoF+frpCJH0A8LmZQtvcAdv8F
jA9eNuRerR5AYNPz+IhS+1ttNO5eoWllYWg6spv8IalKBWKV/hso8KQPP/DLLwzLYXRNxH5Ko3SJ
CzC35oob0i6rYO9FPfxWlB7aJO2FmNf/m3IRZLqW6dazeAD5CmPRdwy6Q9nY8e6Wu+SqT0hJXPE9
T2iCBThLyKJUwNNShHc9N+PPBF03TWqiy/MECf4lrmtc6GhhRKilqxDidiMBA5QgVJ3FIdbnE+RP
fJQ8TqusQlLdY3/l3Iq9pdtVwEmDphqg4yVLr3Ss555jx6ORL0oMz8SojJxWs9cQqntuXgSLQsPZ
hshHzINUg5LZDORk0FU1aH39BzE+NXYkPGNCEhLdjfTvcOJD4FADg2F2CXyTdFFL7JGSmJIy0cvT
DkoTNaBJJmtG0NLrmx9D2MrzZTmhWN4J6H1jXilBRcXk8jqxcHFlk+mSSSpfyr3lyeNR2LXd04dd
4Y1QiSgc8EnUdxSyINWTND1ZJAwk/HER+9Nxg5M/GgSfVAaXvRWBtVAgHdrCXH1zEhOn7RqcSGbM
mSYtJKyyx5kELj048pp8Xnx1JxjykUA7AYJZuEwnGKtRhkYaX8Oidf9idWQRCG0VnlYwYMZQARhM
gGkVt/NJRalzn/SrCLsntdiEAa9koMp26uScmznQEvMburDbv3qvsziNqImYGp2Muz8MaM8Wj6Th
AmPUrFcjd2LoUZfjJV8kdOn3TGDb5kpvENZZN8t03dVq+apQxi7kB7jgo8AasCpbhcsdrFQzOT+Y
Gd8KUh1Y8EjyUv99uHWRsOqHdwAKKcVCbXfbSLfoggrUB6mBOoaLBSoewyGdHOS5FdXXije7NKMz
Dj5eQmzlfJ/YM1hQ/C6OkW/jBPDs1MurnKaCsTC1G4wKAfdHELLbJCa0ff6a31w1zuVrwv3WyGvT
9LK7mh/5GttLrQIRbKGAmdxpfUtt1nbjyu8lijcora/E+/aANPe3cvdMl/QdJ685T2IStRnfojif
1M9lqYcpRZ5ZDChiNrfSUH6ejInNTsrxmSkat6Z8ax/ihQQNnJgKlU1e2g96GizkPmndO2g67obm
J/IUv0Zh5cGCRjoZVCezw2c7dX0qP4kR+bbZfomAVcMj5gqK80U0J7Pqg63a9Ddwxf3TrHVG4pfu
tdEu6N6tw7HsWczy39lizuP/X5wNd82eFCOYUCDiHJLkfwPO9+fh/DWfRRRkOyn4UxbHKoPJ1vbN
xr2ceRmqqmTvbMCmzEu8qvd3p9gSM5birPuaWGuoprQHa2f3nzmQpHE+HO5u3xgpHfh0X6sO08Zr
gJLqSIUY+LJBTuWV1R+pdgaFA+3WytDl7OUut2ZDkBGKxmTgkjV5d+A3h1XbuECpl1QWH+vrQAQL
IValqwm3B4QZ4I/biZwOrI3igTIfwtVh8qNzIe53fuCC2zuhDdmj0JCzU6uFofM4tdN+ADUWzrla
Hqvqk1nHaRByoe/7qQNfHuJyMd7891k9q9/1IG9/apBzdb7sRNbMBGNv9PPwdLOhdOqszPW3uF7U
5dQk6GsBK+hY2iL4nlJIRBxAebpaDtZj6TQXIVktC9pVcjsiDQWpvUAb+FTQz2fkMphHCGGMSiFK
QUHGXJ4lX5e41BckP5RVs/fBF8sOw7+knKYTmX2L+IfR42HOneCbziEjs03qZtNrMyrksstx1NR+
MbwMQgPjumGgvSjLv09krko4UHOXKrjw7wDMJzyX5BNGvQEJ2XHCKsvF57XY1PcBvgLWz4IAfLL7
H+tNOWraqw7Nv0hO9ai8HwMe8ymXATb0UKPgGq+mJteShlvgoJ9kc1NdM0iimy9/JO1NMMaQQ6jJ
yXG5RZsWW0o32Bf5ShM3HfK6xKrZ2m1ALxrMHZN5iCFOVBHo+jlzXvmGrxVKWBJ0fPYq/wugaEI2
tt0EFiyrEJYZdJhXmN7hJsv12R5as5aOkPXxgX5l5Yek5rrBoJ2IMyz/AVBrCLQ5omRN386K10Je
iXkeaRG7LipAuQ/Wt2vgKjNrEXYhJAxFQYxpywo9ZpGxcNMcRgnQQIHZZtVhCTmWPaeNIeC5q2N2
FvcnHm3ELz9v3hEAYP4XE6Geqzvo/FNB6wiJi13c5nF2HAtPlelP0dn6fIeU7QO+HZf9EGfxQ3eL
vBblW/KDVyCWs/envyRWRy8++3JfPM7LacDSyxFqUoTdSfXMSkwNMdYr3Hc3H13fQDbBb0h3W+Hz
n3XQafzm/+KuVr6HiwfsfelbL+Gu98VA4BF2UDmFtwZYZyNyK5RIdAbjClgpNeIDUvv76kmsvblW
KyCf95cwIpUT2imdQYxfF3w9VLwhLI3kSki5TZeRv1e/t56irz2S9UwPaemOmmrdlzj2xKMysJXn
tJabT3zuPDxDW9+qHgFLwc0OdNcmiaxcH1j/Fobq2eqFpQl4uLuQhZ8n3L6BQZ+WkaLrU6OA1cGx
UyFBqySXKB4+a+2d22XSgKYWBq7YazwsyeUTnYm0CH5UXSrgVhcH5SJ/KZEedsOwryfOFfZWKRUx
BF5EGbjDfMZQRzhvtcyqeAgifkkPIMZ5NUovbdEj6jX1pmfQ1WmohOtjogXVgJWfD3sOc7Acsmia
V/O2/0wl91DbjGrTlONtaqGzzozW60pXg06s7QKmCZGfXQfWuQfaQ2aGLG/pMYyoGijWUSXHl2+l
iTMUlwBCWTha6pm/2P9J6qcQWJhksJTC3qNnQGKU1cTvmPmrWsJ2dlq4HsBrJQrNgvQCzf7RJqur
MRC3j4Lw1Vgg9SJ7UBiIyDbp0BhEwOIiuSrNTzFP1jxnmxJ0LntM98l3BcOOUq8xu+qe/C+qSUpC
tnJSSZnU2gOE/wEX0ifEwPYlFN0Zrumg1a1mtOGf9AvEGJ0vyKWlFp/CQ3LcjDOGjMEi3WYvGOO6
+T7oAvTRHM0kgAT7TdnehWncvRLHEAEIFg0pf5KG7giyxlQhHNnx1LEzBsjWO8xylzp0l5IDDTVJ
4B74E5bzjUOI3rfd043h7ZqQWeax+QP7Jk0s/X4gRXNcea5kxuSktHhL3IA28B4n1ZQ7LaugTDjs
EBeNcj5ZAMVTgXj1Bmr77+QVk/9GRZCg/p/uhmrd7fSXam5BDRIpltlEGSyYqYchMGZ+zvZfJPSY
nLvZApCK3Etb6UYzqPg4kd3PEkOKgRf7BFke98PacQkjGirML13Ed8huEeG1DpFx94uipcFGhqT7
ou0a6oFEHuumyBdyInx7Nx51BygUfHfKB9HMIJsz+iwmEKtVV+6/0sq4yWQ/QUrEobLBUrLYhDeA
a2I8irRZ4Uez4+/KLb9F5K+5KbxgCcavPgwxkdqOpSy5xm/t8rNcghU2eNWgAXSCr2H2iipFg+Pu
sPmv4PBAL4oJNt2IYqedE9G9cbmEu4GwC1IV6A7Ji8KmU0NtjaA/jHVwpuYqdqcKtMa+y+NnwVE1
LEc9t8vwQUYOazQpXszsZNJKOGwJoxdqa/GT3TzBv4AR2OtnjfOaMdUCsRGxTSnGZTG34I/4ZooA
bDc5rpN2hNQvlvvxj/mbGjdO4nNVgZ2CvT1mEcJolyPAngAO8hmvlNZngkyXU/VbwW4ZTb817r90
V36g8JmZ+Tm1m1dXbjqhqOPoOdkuHQrJfFqfchkbF5s5gqY7C/iftEfsgY3nmc/lHD1naTdMVVUi
p6qZfI2Vjb5+4FXxH4na8sQ36Glm1S0YGvD4s6PxPmDk4lu4Xq6De2nsyKzS6yfOoJQ4neX21liR
8ooaiAAwBEmTwL2r3kIFWKpAcvWwmt4YI0LWwcnEvfj+F7Z3+MHMyJHB10KRRGHSKI5jXfOj9Gm4
rEDQJvL2+u3AZ/DpUYHWyBeckUGCUXNSs1in/QUcR9sulctOvo9iuwPvId08cnRPTB0neB0GxrKx
lde7cVra7fO1KOaqZGFmo5/jTgpF0KU4Ou/+3c8ycSSYvupXaiFIwR0JQp44A7hHZGyprFHZOZcT
44/Ae8CLXWpBJ0T1GEfTwnpTYKc7gKmkJTlBmuH7C6NymW+JJEdvxHXvRi6Pq7yKiOYFpmy3LVcE
P9imb+RMHfwpZLLyWOncn8GlLTV/6XUJGSo6cBHaJh/qEoOH05SANujkIPuA0/U0v4NhlDnPRadr
7w8zpfRNdp9mFRhI61Yit+GhRLwlq2enDrYKJC9QjD/5uVRVfPGI0euD9tL/r+0JK3ils+lwpQm0
lUyfJQrFtG9BpQXjuReO3RhkU/u46f9Xxb2AHNxHSemhLaSuSw7xMcBj5JzX6qotl3dgdVtNrsPK
oFsICJ2Xibn25Tk+qjbmxp3T9lzfxC8Bb/K/MHrlI3TDmaOrTdoQtPXGJ+CB+hyKWBlkH0Xgdj6U
rUWpjBOL5YahX09tu4Rl7qu20WZobMyxsu0LgArDpcNmz1hvfCOAX9vLskU3303NnC+zmBK3YILU
ANm/Lnhsmxm5KV0TnUGx5BpZPCZw6A5sSXJxfjehfixerM7znroNINquXQavBJ6iXDejuTYBoZ9I
ASQxBp4nRWMxaEJhsmyL5Ll2n0eLlrjW/QId4bNUgcuucakO4T4r55iNBfdN65sHrFUiTWjhdcI7
UHWkUXwN6D5UyIva1pPFv0u33sJJIYP7piAbCFblu2z8IB9FX+4B6fwc16hJuZGS76F549u2COQx
N7l60uyZS8dOaO93TUK7gjkrOcjWCvMXqw4rImBnGaS8UI4bkpNGMBIi7irkTRiYT1XApIsE4ESI
mP9EE116DeYPI9FBFXFS3yIax5Wt4auOnw4o0TScEJOhPTP2Gww0dLJk1wrLhRZ55lynNG7FlO9p
pyFMC/rqr/xllsDiLigzoXnXUsewoC6kSDxxLpHmeHDOAeBUUpiYS8kkxlcjHdlgHZwLYaFrH7RW
NZoGLvLlHZgr52cpEV75dMLsOjugiux2JJNQE7k1CIkN5Mj9vw8jXZ+Vk7l4Sbj7llNKWPmzgkId
gB8H/VzYHha0bTBERVbcvBHeHlLxzrDmEYdjX0c0nnBmIj056bBStwppLE6O+egeAcrs8MWltgdu
D2oGiXy0zVMHh5npRseIpZx1sns03tsdV7P0SXM7hSixOVBSD/ae5fWf1jEVQ5qIYUarHXXW+MfB
/MvzCYR2L3CuTfKrxuTrr02SJo8QF56x7/Y3FWTwG8p9EVblajKCfWfvYNmlkolfkuk8YYMLTM9A
k5pWAZobu7mOH3awVUEa39/t8YvG+li+dhLnB2CD0SjE3B2SBvgWgHtSrrnXsiCMpo1hqxEVKUGG
iFFdbU2WD3XPBafHpIEPjPqbSSorzOcm1ozzP4vWXOtnQ05gFCr52RuzXlM0jhxdHTxMO7CO1FN4
IdSgnBfHtMlKmgmG2ZBEGujlEmPbMuVBSTeiGCm/YpHIVb5S+bHwEjDU/N/V+RG9DWuBYkQ3pVkc
/5EpKEDCNPTs9Nf28/JW5w6QFbV9nheKxf4OaAAyNqJ85aifKM4ssff34FajfsEZw1eYC2RMpcBC
goPXg6SrgBx6dRwQ4LiPWB+zSWN7k61jGokvDMSqfN+E9j38btcNCMLuhgpk2Xo4lF38v65DO5J/
CAGcL5+hxtbJ0hNf0FHwJEy97yYRG66VqIK/R/+7oD1fukY2h1h44jY5qBq5bWvnURr1rU8Fav+F
lBGL2xZTd60hVqdWVFYXF0lckb8XATrezMw8MRDmC+qJl0lQ7ZQjPT+TE0RtniKmtWVUflp64rnF
awBfE+lt5FaAV7eAPZvixflvl1Y+tyVejNVGd47jC72DdyaXMTI1D6lrGh+q/J68JXWC9kIYZLR+
vG8sPqNP/h099nzIC4pPWVH4XPYZBRMqaYxcttsvODjbR+4FAeDGYUymALCVu2JnJ/1EqtlqXpCu
MBkjhQjdjTdLK+sqy5djolSIZ9Rhqv44fPvahnXbVPZFcbbsbDE2G2/EZxYxKmbCSFElkJLYR6db
zlJIZLvJP6CA+1vUFDC+6ragt9EID2REtzQEafAaKCZ/9YrIpiqqML+IYLjrtyEPi+vPkFHQNk+w
pNdRQUPLiHT/o7E7ZwbK9N4GOrsReyJvFdRrLsWhMm4X+VWlq6Sw48ntKZDczKS2MawXTvENTIze
VQN1mOYeAenOLtDa6PDqoENiyclKV3iLggxp6ChLDpu6g8WJv+VNAxjwa8HyunHkHWRb+qzlxKWS
gqeQsbLkN9W85PxcMJDJrt9aRDBxeRUbmBYB0bjBS1pEG2/iM9k1h3QwHsXsCYV94kO3cbZcCiGB
uaXp8vORIjT70eB1EPEekRkXJMRbp1cwcPUdD3M5LnAA7ukXftyHwMWLceZwNNeRAc52GIQdDzBW
cWdSNYloQsll5Ux+2bdlSvo6dWNNatUBbVMVXSM4Te0M/DkRJJ8xKGJd2i8xfLSKLrTjeSql/dII
FRWkOgn+O5k4WCl2ZtV7fD9oQX54JMCXNTUigPnLK1mqhzGDxLI1bI4kkETTxYGqdyp9GgOmDE5L
TJqN8FkqfWZa5IaN7IIbc0eCCBcXZjj9AOt5AraEinyDmmnDP2HjaUVIpY3ORhtIbCARNab0mbEa
Q5M4NTbMc08kPANGOEvfny8j4ZTKEu6ua811rZYddriHUlsnD3b1b1yTiZxtidHRm83cUBbZi2vn
qABuWnjtG9CnJZfCm8ss9as6/8qotrvwjckcjP2NicWOfVXDMg5esYEzogH9VLAJdY/8vkxEh9TZ
vJeRhqcF2ojnVJuNAGsThk7WN+ZrJ0Hi0P7ajSoNAMCd6hnFOKTujr0saYfLAc1sddkXYKnOKQRY
0inLsV1V09eyCkHqKw2vV9g/0OBJ4rmJEJK5icEgumKs3YciKaN4a/mNeDl1ZPchFOe6L9ORCRiA
j5bO09s4ZuFCjRQJaW2BmCBQr9ujQqfCuTpCk8dcxqAKl5u2HvEubgE342ieXjrkoD8nHg/KLF8o
bXNjiAu9K4wSMg9w+FjOjJ0scFOXi6wUNl7hguFxhnxGIl5sMOoFIqCpLHRcvL7r41H0iRw6Gac9
wUTyJIfzAs9bsT1cpn1Ugg3t0/Nt01T7ihXGBkUIjA8Q651ooVstB1+nPrE2rdAg53Wi/bfVCyue
Dcxh16VMy4cfSVGzIrSeMxfAHx4WhNAoX++XvRHaTzFptNA40TdRY9+BOlHuDd2WcV62nP134Mkr
0WHxS7lxEtyaxv0PtiO8BGBvNRCql8du0vPJG979fEIV0QJpJGUFAm1vTpNvBB9nK+htIZExjtLA
P0nXGqAU60vsFcFp4C899M4RnpsJdaFcqYwrSe7UecrJQqkyq+MkYNyVdUEcwzlp1npODOqx7RH2
YdHfelqNrOBciXrEQg5RYbt8bCfaJPMKkCUlzmKD3FfTuIGCM8REHF6vzNJmhVS3GK+s6GWqyf9d
B1UC+pzEsx7bnVvSe04Fzp1Q3OnohYn/buKD0tdJ8Y6eJkNXvp1Enksv8tp1xdfouThHBDNoP7d9
PhHmhOfr/1A4EulwOPoHUeN0WQbRW7kSMK2XmhP/slSLre8o0zIMOUAAUjdDvDB0xEsEeSojqVFm
Bgg8PJ+aFb8jSTMbW7wOwqKKdUQG+6bb9MqvZNoFZF01JE6sy/zkPS9l9XoDP19Py+DwhUuIWEVP
Qyf6imfC2dnznjTIAkuvPizRgj9TtEE7Ff99eXcaGJryFZkV2zrzxXkGxgA1XibnGTRXrKl2u7WS
+L7kxg4kbR4BfkcnGyDIQcmQyKhbmIsGIbk3bt8kajGXUcU38Rz0oDK2B3KmN+i7WtzOQlAeLXkL
fP9vxODQ3rqAXl3VUyFicbocKDyl2hfSOK8ptfN4CLLSppQGG0sDiEZJZgOG740zBafECpVWamLp
g0yA67PrNmiyU/SoPwewGPK0FdAbQ934VK5BytUZMriEf/g/Zfr08smNIv7A8/oH0qJyiZBnjBwq
+35sEQJ/ZbjOBWGYfmqm3JKmbBt/sKx41zDiwjJvGBp0xl8B1WQWNCaj/AkJGY6sZibQC8MGOY64
35AhP+2/UuwFHHECYAOrcHER2q/oqiX9UFYdnUjt9eaqmWZWo8EedkK1HJkVNurQnyHYYiNsrzOL
9dk7gLPawJzduoqdzLNZ1BxmdfkXyv7xVZ7obYgp5u8Vf5etvhz6+IWKT/IjiY+WRJlb2a9tEmjD
1almL8SPfe77W/SKbpGx8QFFD4sP/ygjFvwVfn71VQJQnAYYOkJ2vY9jKYw3RZ8avxVvqXLHiVSH
PxXNsYYLe+n0paqE/8A4EmBSWJJ/f2MMiq0yrdHb3WVvaHSCquHJxXeBnS/b0k0OiLKFmA8GvTBO
LTVSVrb9Oza9wipmmk2uEAaYandlL0bL3qcahSS1eNrPKIaYPIxCX4IYV6gCC6q9xGteRczuJ61K
B8X7jTDnAgD936fgCbaERmiTbzJ3lxeRnoGCzEIyEz7jUN+TOQSELqL1AbOAljGg0ESh3DA/6XGA
ayXn2bsCn/a/j8CvMAM70VqyGgH9396JQJ9m3GYWfItmiOOw0bi/5aKL8xWDn5IPdqHmfYVBWHGe
0XUjnLXVpycYs8m1t4vl3husrKC2xMjzMm+XNTRehFwdTa1YROGxRbdXQwkZphMimEQ2I+XlSni6
Kg/2Oz74dhY89+gHk2ReEMfXqMXppafM5NfeV0KpqEf2DlRhi0ypm3U/5VrARIFrOgdMHGuUyzkY
VYvSrNEcLtLb49Hv23LmdI49YndbtmPOBpyE9rHCNvaQ2du5RaXDsw0bblT+ABQy4dh5rvvC4MQV
0NAjH8c7F0OrKUVqRvz5jucgt7vQ5Z01fZndLmvDuule6JttNqfMZoCpDnRuWX+AW6meGJniXKA8
s0zp7MgL8TCEUL+by04LCX7IFDuGFiNu8XrxY5Lg57W2YfdFgwwGL5oLut3+z+toy5Jj8hPLCTWa
Aw9axbin7/y1v5qTTDlN3IN9vrWiPJOJHAEmNmM3B/3mDmPg0xgfEjK8xXhiRfOo6WwHajTvHV81
4H/k+ugUXfrzu9PpRgXw90aKLLn7bY+zIwQSaWaecMJJPiLKRG7r/60MX7NVo0AD3sZWIry1eVqs
Up6fuRjlYUfLF+6V2Q4ih5PYmibp2aqe9l1THQIjjFsnE1XlkMm41vRZz2QIfx2peLifPnxCvOc6
MiZj2fXICPPdpuZXF+sfKC7JsqlZisLxXxDcr8VZ0uOPcVoU4Y0Zv1Q7v/zLTy0VkahaiV7bsLJL
XrTnMzUtyF9AiXnoKhCQzcHVd5Mh2FnWXZMnSHWHGBgbdmml/U2gSNFVP7x4XwFjNoy5rCn05zEt
pPFJ1hLRNPboeeAw27wkJMVUa7bvcfOeYiD86Q5neYbP/oltd/I9ERhwwfT6WGBM4BSWLyWs9r6t
p1ULGCqayW6dmMaxUwtbHWjexfm4DR18l5ldP/rV5mEYCcB6JT+XzZpAO+rWOOHlOLUHGoEDRQ4q
3vj70xzxtYkgl4AlqLPZaHWI5tmqGrb6hev5H9vyvVmOcR5zep5y36qTqdeg2Z/sJjX1QkU/5j9H
NHpcvsNVSdMGDQl6neXZkADLsDpRYNyxNhYYAf6EEXxTEQQzuO2sd3wePkB93+wh/5IcYB5lb+He
6myJ+6RBtTiSV8HhIPfSFcGJAbYdszZ80ozhRslqdelgyxsm5tM++4D6cbsClVRV2a2FQfPTi2uG
WNQIvab06O5sxGGB0JsGgxjFleSmCCw8dczzvIxYcoIOp7TqrWylP0dwQ3rDUt0uwUtt5hVwv8Ru
GIymeTDt595TKb05HIcSmTnjJgzc/C7qgMTZBIaoXvASaHGXIdAmSNBEn1/S36Zr7hLPR4w1UedW
AQnf1ZO6Og7k0+LRv6Qy9IkpXny2yQ6loaTFBrGmzv73OHV5oAowUTCD+QIkCFQyC7wfu/l47aIi
yDv8cXgkbaQoLj7arI8HL1g3oeAvCK32g7N+9gFtG3FNXoUP/R1AzJ5pBUJ3WSRoKueJ+/wHombd
WPRHePVOBuFavFoogOIT9A2Ia1X28vojounoaGuTqk+1MLNkf7+tqXn1YED4bFDyjnVq9K0GbfzI
2So21LIWlP6IaOF6eHQny1ZDr6dG0xoL9rVJ4RlxpSiYM9SKoqHxza/ggcHdRLM9s/4Yg+4staPs
0XJMqPShHE2Fy2nUF3cd2ObA8UdBCmXvJ3svTqPALFdEXO3g9LDhRcxFotA7PAWGrCX41HCxhkCO
vnV1ANphdBOxP1Cw8pA81rV5v1+UkzMPhcxJ0kz3Q0+70R0u9lqL1rWOoOVbL76Eu0XESrS6Pmch
6DygJMRmFR82g7WDhLNPelW5ri8xbVP8wlme1lHLUz1GL8NRf1HmYTYdeVghEc05mzXODjO6FHV/
gW4HIjggmwy7vz1Np6/upV5ppgihCBuj9sG0uLG19Oc8XVa10nPiC8ooZE0XbQBsNQ6jmMoaZgaj
1S95hDagE5QHPNrrzy6Wi5TvM7SPAS/h2s1UGTY6cqcXZHfLse4h78OHQIZXhFD9lO0T34VuRqSY
J1UNYiVO65maFiDhJaRQSmTkDPXvgCn9Ww4K6Tr3VGALuZjmn31blu2lYvM8Ie8kaUeQJGqgdIAy
DN9bdi9Wym+9BbMSyD/a+f4VHW//l00D0eKcCYBtEc2RI9eUQMMlgdQA9F1rHQ6VVDRj2Kb/H+ip
ZoUG98Z9dSMbLUWHTRSQS0Rp3oC7dyOs9ZVWZPZSFY0GNytKoPO58aAnyUoaQPXKe2ZkJW5YRATr
XvCqa5uQgNeQrpc5exaJLNiApvMuCySq+FVrCFPbVvV4Tm+4KFHBvQAIaBfZtYh7dds+y3fe1ydj
LHWzO07gRxik+1nDHCg/jyd7necx454yHS1H+ncr4ZXLnjo/psdg2XYS+Dx4VHJCrRbAp5aHGT3j
2CDfdfw4TxMPqtNj2QxGVNZ5hhMeCe3aLZvczH7QMS4N2wGQN+oQrOdQEGx3jvQnk7ZkUVOYq8Jm
JJO8ISSEVQyj98iaiyCXqOCU/1VJIsxW2tKxncORQpMgniprMSe/U/EYnF7STceGabzMMKiUa/3l
dVXqfWkZjHc1pocvJ/3YLZKEG7ix/nob5KVi7g9pbKrl6arc8cq5Ae3bpeYcRoXVqitbrSPTa000
QfQMcr33as6/F+CwMo8BdVh2oJ/OL+WgmT9LQVEFbDRBpkvEGtLoDdY9s3XvSku1JSBQg+er1zoG
uQccvFvLjuaN2dgPPQpmMeoq1GJHDtRLURFwifWHJ2E6C6yNeArCGHuqp5S7jyhuMCHK9ilM4PE9
BCYs0/e+UAHdlu30bPnf2I+F8sXhuQup1AENSPgsEZfE851WiJjy8Lmh5T33mpGv0kt1Vbw6uvMP
oNjFUdDLPZzLI+vsn0HxCUznuDPldGohUhFXniW6vE3My0GiyOhJ8K1T87aKaUTCfsIXZ8BluUGq
K2bDTpo+0vQZzez8kQjMQk+jPYN/5yzVzZHfdg48Ph31OV0fWsvdoFx6cQlWCQ5ub8hrsHv45z2S
trWZzYbRUyYfkn05JeYJhH0aOdwft1OcH/ZC91zL2WjJmuh1m3hz416ZLCsIcoh88rDGH1KX6U0+
pNXZD2ez87Nfh4hp7E+ukYuCpB/THZLWIRmm5R2ceoSkM0jMbdwMSQ8oesSXv1k9Yl1ERDH2GXNI
9NXpB5rKmEgRfI+4dehHi1K7OtROV1wC2BBbukk8teeFgSOg4NLjswgtvy5YTywEGWJeNeG7164T
BeHbk+Vnr8f9nqWh3TCvtDOqHtrDBp23tvOjunwE1/4H/RwZaTAEUd02qBbdX2mMoBwYQC2lrC66
Yf6AaO0jcddsPGi+CG6E/RpyPg+RO30EZdauU+1ss7xgPHrfKeBMGc3GxEGHNXANgwMzWDkkQJgO
XrbJoKoQMlO56i5m+ZbVUEZ4kA2zZ6e0+tecOQII/B3nA4sILm81m8yC5nwwlJP76VFynue0PJbw
Zllt3sesgQOnfoHD+whBmwnTuJetfnR3K06aPQfMJiGAW24X2inh8AkQLOGGNWtk9kSMh+qlpdww
BX89MtjTbW1gLiD1TjcqezDEkZYNh9ReF/UP6Zd6K52aorsJ1IdF4qLdLmK2CUoZ9qSQ4ZUnYjo4
IozlCNkIfC3beG29XmkKjZjvSpfTJn+RH+cw9+ZlEnL2B/OXTqbhMyIAzZYPDIyf3GZq4WlUHgkV
7BmhoN726UbAdWcpmyEKv09lj8pYfdUhHq9+nqr+OLLZTcAy44mQb+luQ2Ky9vR95AdhPlqBWjqs
bwz1jikMyo00QMjjLtcgp9kSKfAeq6I1KrkM4HhSGUuL/uU8CwjicXZ4IH+4XUoeevglklMprPqs
vOG8XD8kb8goasDPX0ON6t4xrwy8x/vqcCjb0YZ5RU+uphb/vz5w3tKDscv7nPy2Erase21APHLO
JwfcKfDVibKa9lZFK1pj8sT8gmRKQXeJnDo3FVMd5/BIYHETpBzYNsDHP8t/spDX+QSd3Dz/zNce
prqklVQqM0Jw20c8Aeqw2bvt0NuRt0t52TWy7LcW1tWGvVDQJ+MciDK9Dem+PaQ4x9mrYpoMrCXi
8OqXl7QgF4X4wjjg+eGgK4WHCWMYNzPAhPc9sTyRVQXHm5eLSktwL49tMs6IzXCYvFDusGWwmF5t
tJlkN/1DGsu+ouK9kijfuOKCWsKmWwXLyasY7YH6ViRO7/dnM0Px8TPRHsVsCxlVnbmZ8eLCcki1
WwPsVmjG9lh+m5/Fejkov5J468AyAa5KUPmXT5DhNNLk1LZixR9ynb6hts8IStiBipx9MihURNgw
9hfH/gox/BMOe6hs0C8XCNqauh2TO/W6QumHoJZ3/PtjRTYOT3VCEAM10F25nC3+6i6k3EQwmFhc
apNf5ff7XVXsZiH1KmkU8ljgNMA8+i8wyjLBeRAUAtZGTFpaDx83whi7OsImhPACuvG0A2GFBmVj
qyLN/C7htBa4LypAKCbHUnTaPDyItU4d4zVqaANt88v/nljSiayjjALTLXNRwDEj2/k0xW4y/AEi
YbKvG2c8bDxLdnICBVTKya03mm4LzPQmjiVpj4PF9NLCB6c+qdraM72NIiKjB/ibBjTs4oUgw/BB
qmYfirM9P/UjyP8O8DqI1681CJ4/uPrkxwVCESAU6VNAXT0w+nJgmgBHwJSXJ3DpPsu7pGpgNbpB
8e6YN376OoxKAB0Z/Sqs8m0H3Ew4PJnYOz5L8p5H/zeFz0mrRrX1UZ3Y5htOIW07lb4MDupU4DDZ
5dQtk2Ey13ZZFWUsEZIFrJcRyr22cScJ+1rqZVg6G1yyDp0fJq0p7T6Z6695QmQTbFA4qDNPCvpi
DegpeIwSHkFgXtSpEGrq9WiVK7GKIhaPf30oD/nQGOcoP/EhFrn0OTKrHQNGud/uXQlmepBmBnMo
Z7uOf/LqWsb9Iw6rPKgvMYliJYmWQyBiVUPgw9CYHX5bUR3HucbLRfeZpwwkIFAdEuKlQdi6spVF
W/LL2brHcl/MBmJmSEYaz3xHw9Lvqz4rxKM852B57cbgay0ypTfZfG6Oftp7WzxNA9H86tJMaEY+
eBL5VhSP0ooJyE38AX9KNaoWeSHdDyBt5dgb1AQukzBgIZT0NbZl6nuUhSjko+dOQHp8fau5gTCY
rQv5piGAiCrENVoosjwZR49eAWYPscB34x3ChGh/ffx7yjkgzn7SUrAWnoazf1eBQq3lZFBD6I6j
lTs3gU7X6zr5rL1ctUgdWXq/5dNss3ozKtZiz8H54gB87n2blTOPTfTpGx3OiwZqtNChlIHoGcBw
Fqs5t6ndXovWWpOZ65MLYUl3LVUOMsiI+IJPQE5mE+elGabsRXzfroxmmh08sPndWDUD+yKnLLgG
DG+FOqDvV00L0cZ0K0igDGL6vfVdJEefueNnMhkwPC16piVx+xoyf7ifU3vaMmkvy/HF/SiYQs7t
+XgOrwj0S/SiyFU19jofCL4WuCwc1cI/pC61ds6xFvh2AmU7YYMYGNEu7gQGrF9A0iXbzOtwxYqr
KVzFf7b5OzRJ8t2wNGrU7gO4bu/ZP5+zZCdLVdqWanSZ8DUnz/zVyxv2bcjXdVQ0RPfNS+1Bnr3I
5v7MtR7ErDh3BodjGztQthb/p6TNrsyKjHMvSL5CDFGvN+4sWtGYeUFx/4wXeZrLsH2dnWIEM1Nn
bfBuLfm+xuEeuUkPj6MPnx/34BuarXSv3cnkTusUroaM7g7jWhCj55CNOGQNmi9AtVr716iirNke
C3QDKrPF3UVmn++vtJHkRzvd9MEVtg5elNfk19tjESO7F+od6m4sT+OXREEuRvdD+0IN45VIixsV
DODAg5cJzH1FiKmdDohqdhr0Gq3mNVBVP1/n947OpgXAppymmcv9qXV26PWpJ4u0Gr7xxItZ/yf7
a54jRXDGaRpdOeqI2XUJbjfvs/8vF3NCejjjy6rEr/lOpHeMt5XOJFqKc/Y4Hiy/LaLVLc+HxdbA
03aIf6RQu2rGeLS3t2vy2/NqiOidV23xbr2oatSwdOUcijhRCF3t1lsrAk4wJRJiQDI+bINxEEVu
9zo9mP/Nyg/0C0DSIFfo1A2uTk+EswuCqYm3UR1SGrvLhmyQnWUrUDIsvtHfqetZgbkgqZvBqy9A
5FYF+GmOwEOspuJRwcCtQaFuqCSR1dBNZtj8wI6UECvctkzRfY0D4fXWG4tleS3PIGM8t98ZCvn9
ZVzzdiw3Tt3785nOGyQMx9abySC30Kwg1MGqweuZGzJN4WAgeO96OfLu8EEENzA9cNbPJpXAh8Uh
Bdwx41Oi53XnmYP9QCyjQlXQ4D0CFFI4zM7OoPnWdpIY8sXjncUFeQnKu47zqq5fxEwNRNMoHkNK
E+BbEgkISHoQXhfvOxK6m4Qc0d/7z/K/YxOlT9w9sOTuQmSjjm2PTyl2rvcxHkYoAjwPfM3+ShKc
TBgh+UYMOzNlsIF30L74bOf42HZz4vuuuHxBNBFfTb3EnPPLkAzqWaYiP7zjXznQR/3Mc1WDwVtc
wpp4h7cT5WQK5DyIaoVzQARQc5uS3rkAFo9cmwJ8JI9CWFogJcmQ0KMxMbrz0WxZFgwcYYQqjaFc
zSwlED6cCrkxxoYFpOntxG+GfqNYImz7mxb09rfYa2DFhF1LrhC2mAoQjSAp6yaOEYId1aErjUj9
E1Vh8H5/+K6WHQwk7Ibg8ICRbUdU4vX8+OWm7DtvLrE3cP4mWxshFVSNRMR8txDSAhilnNa+i2w6
tSiSEZzHc0C03upq69jR6rLHoAguh/GYUiXg5zlz+u1s5JUCWlUuEMoyr1PRsU4HQLvxCSeRypLP
V/F7db3qk+fKdPICRU6rrunFelYQUMrNGRpZusSYgGb9b2D39eO5X2Svv6O+MRGe8Azfamz3kBMq
t00iibKwuJKiA9xK+VfUg5Q7ID0djoIb1+oJ6Z+zu7kjd7esN4mryikfYDsylISrD/EUf882HvYy
HSOfVMp8AZMiUxgwuYmUNgPhpvX9xgTk7Hu6IAw1xMi4OyimlpGFrLK5O0ZR3LwUsGW7XsNnzf2R
rZvoica4QjUqgQkJbjWCMayaW5N74ElPIvTjEF9HbAKR0Kyohi5CFX3tSbhCCuhu3XkvvaJTRHFp
48rJ3jaGrkPXmavfVE8ZN+FIJR3bAznsGZXejga+P56bB1oKkJNsxPn814F+WgBWxLj+CilWH1N8
e1ivS307tZ03InZZ/mkhtE4OQEtwseTjH94Usv6DkoV+fY20JQYqNbTniYHMX8zyu/3Apr6XLye2
sPD980aPo479PI4/z+4dg6cM6L6HhXevvqQeVwNWYt7kgonPmEZ65t8eh5S8CLsS7fOJA/qlq6/S
qs6ZFnoch0a43qJCXmWMW+s/2bkzbBCV5982xtg65IC+MLyC89v7veb98p82whffCT3V61ukoYYC
J7mMIz9azXQl5kI59Pw/DxzZnklyOGxw6PtM1klcb4jV/vo8v7ETEf3lqH22+6fZ7rnWR6oGzN+x
jwo9skfMP1DMn/tNTVdd2beFUcvc2lU2vEa//dQxV9pB7Nv4uhKxHmKXGDPOmgGPNOSXx4SSX3M3
u04nR0IXU8sq/zj5/w2IecxlziXyzg0FIq+fxlmAkBXmbD1uAHrhec07Rb6FEOg/zoe3ELZHHDgN
AGlgKTTlHjem6p+2WCAdKDtwlGs7aytg/nAxbPSHqO6jSZrSbHWmPFNs90E0H92mIgexoY0xMCaq
NCWY26V9vhWXxJs8IihqvAspzY9XKCIZPy9+eO8z8NZIB3l7x16vv23sADkYuaFlhSKAqRT8q+Tg
biizimaKUtM94lrsJceMOewk4mpYzj6KZqM2oLKZLIyyELtYdpLrLw36WjUJXhLCczNftPCageEH
G3/QSkd0mo5mp+kGL3tAhjp1LG3umqQhCOWdArQo7sjCBRBdR2D2h8U++bOTrb2gfA+P0hjeSNZE
QAxbaNa5YZs4cBQ1RngpKOoQRpLN1542RP4VEuKnA9kIgPEF7u8y7tNgsvfsrrDCu4OfNPoCxXsn
d70yiWqsQ4x+VDvIY5zk1xv5qv8Lz0OajgupF/+23vDLT0X4tt7f4FZa2ukatxSGvYmCeJMoHfme
5eA9CCS7OixHoFbcbkMlcOisNaZcBRqUEERr8lNaoEBbvUnfUBTRT71kDx+zUHyun3zUVCTT6vVE
4bbZTJpI40HCJ20poWCQXro1UeQQVZ1DoO8rxSV9IBOc7Uskx8jjKpdQOcmDT4nBelT/NWceF6j2
DYBw5r+sXUvrEG3Y6y5YNapc2BXCK34JjaP9GmyDGs1ZcGwy6KFAleQTopNpKY3ilNt5z86XeDaE
p+4AcCwlJ9u21aT6wn3HCPANEhITD6SZEVXAqNKmlSXo7DDsl109sZpGv9v+ZFcdZ7+y5/qBiBT+
LcTD8qs88XhcKSdjuPDJolcnuzKkklPVB9WTRRpEXhTf9sXcJwvqLeCLX8i7t2LcI47Hnwfs0XH+
WdMEuOWvaw/hlsy1bWazCnj52SQjPnJ7S65E87WEzOlXwL0YgnSbeCwL6H2Li0jze+dtiFbd4QO0
E/90OUFxvhfZMFs5d4JuDkhiuZo0GWOLBMgY1cNx8wzWk5dDWGIDUZ1RMkpS8TM/xfZuLJcCfLfy
xy7cMbdmCJtM8R/4PlT/+pSk4nCOXl7FZs3kpck3gIjAPpPC7ASrOMIyKcTTEDri+SE+Gtvc7g/C
eBzt3VsvhyH1F5CIJ0UZH7BhhoizUGf1ZhpB4vXIO0DJazRf5jkukv096TU3G5cjXb+M/fQfmyip
6MZ+RCdsQR8RWHL5h2LDW/IUHG5z0/Ttof8cSzt6W0kHY+YRGF1TEvTAun8WCN+RNSdZqAfDOMex
97x2TtoJ22lNIRA/6BfC+kWYnKx/rZ0LUqOSe0nShTZuc6K9+X3/kY7LDrW+SSLh61l1ab7QxUID
PmZi0Md6EjUa2TAeXa4LjUvWS2w5J3IOJHfMIKP0ui1147rquod/SEGZ7hwWEkpukmN7+YEWNvZi
kfaVtLWUJY6OZurdIhynk5yHnML+3XvGWKU3uUmARLhvbIL7fdle0nGJTfdZ6qxtUU0RgaHeFsND
r/wE542JLshMYqiw8/ShyHu/8X2l6ngCfRHjR5MyUEMntDAVHSN6tn3YFun2IUaQa+MiaURy+OXD
zIqvERaca6OloRLpq1i+ee1XgMopPpGPQqdI34YaGqdH179Cmv3K7PLvjTBe3xY/Hn2u2l5AixRW
CsTMshiuT2VKmd+onmDT/KXPgKEtBxn8j+4xhjEdYQyk23XDvm3YlZZvI1qTRKtjcP3T5g6YYIg0
xYc0JIz5TL2y1UPU+rd3vWrSKxNJlUv7fL0R7ZHl5MRtO0kgmDGtJOgKajlcE/TbNW5VwZevhiGC
o0jUDe1xZGWcwm+ORd7JPzbZbgBPm+4NYxGSAaM3tQFGzNkJJVQfMmi1Lf4Qij4K2k0io4kjEhqa
ZWiqOTF7jYUvidxYMa48nZMH46i4JSVf/VCs93n2P13L1nUo/BUCEBz/md+tOy3D3b1nfZwvnrHq
h7CdR0LGY4J4bM9g3ps2RxmFnj554DtKGw/v2jRcxWWjljVOEq0WkoOnlJTTeTbuQsEp80nN6+Al
GSeeLtSJG5sij3+fXsFqdzlxfa0k24frNXvr+CoPxt2/Z6t4SGx+sZSmxVjj0eZbX2HtCzyFm+OK
V+tl8YcIw5g8LbnzN9keB4EnMkEoi6NcD8rLhnYUzR8JlPppYQDVJsVLdd9/TIkzGC9CwTFC8QeB
nEonRdhcwtELmsgttZ84yhMW/y+yBRq5nd4Ok2GTmig9i1W7BrxNBL1b7yGL9CzpKH/8RLXk4oKX
eXs+woLwaIqyhMO/dfmYnebAr1rGKgeiiiNr9dTekhQo7NjSj44LBtodil8NdUZcKhL8Yv8oY47x
K75uRxZqMb/AXcqWk+i+m6eJWMUNMVO6ghHpkWDRb8Lso1V1ZaWzuHOXqjZbE+k8hA6G7xvF7F6U
srCEplt893JoUf/VEVV86ptiTNrDrUmiTQe4yYLEOp+8w0xjiquK9mjW9kDGQQJ+5bOVcLWRcXtx
DegTZHEyN258rwK3MvMLcWb2wmh5QpdvuExsjvCeM2lAQHRDFZc7rpeY+qaClxxxiRN1tFU1eE2h
ZufjtaebO03k9cXlll4RY3fPuEPgYJqkiWusCaFvEBzv3TeENbv96pZ16CoaHUpkr0k4/1s8XFBM
c1YT2tIWA42+NVpSLAw5NK3BJ7VM1gc6kH8neqsahcl6QKw5hXp6BUAsUdZtRRzJBs/u0h7sHnnU
Gz6loFDZaoPnhQAOpE74EnIi7w526ojVACdHX3V9hglwcVdEKsgpzwdD2Gum8a3xQsl4q1U2/6No
dU+voy45Gtxr8JHJDQ5shWfSP3Ph2RqUkZ8tMdVumTtsVRxUzGD2FNgy62/SJH9cjD9JRWPDDvGh
KuR1epbcuEKBAFcUnf4gnRSVRx6/agw086BVMk2nQXf3zWc8mzs1/nGamGQY0R/6aE8Rhvn7LZ7/
gC7XAxeiEKp7Heo8xv8j0tp4bt3PcnDMq5zo66fvqr2zamtiZsrcYoSySP3BXzdxu1q8HDhdpDbC
4L2fuYmGkNuO9xhIVWeUQP0midl4fLn7X/hVSfJjkcYtNzQBxLzt9ZqQR2K0H+L5cPRFrF8egthy
oT5qAfpKP2sgPP0RRmoi/1/yDp/K7GfVuLtUa3IQOHXAV9DEk9AJzRnvebawtZJDswIvs5nBe9ST
ycZiLv7l4Co5+wIXCqR8UWGfhPkneglLQlQAJ+AU4FJ+KbgUY9NyxmFpUiE8TWRTTLN+GpZqJFPA
1YRzteuz9bkzQ7vR8c3U7wBhbMAevsVsKhDAspYL2Suz6c4/Fx25V6ezliIggEJYcfRJq5FssxRi
TK8x3FzqkbF8lqO0b0rhCrN4FRq9SRTgC6V/YTMmpLPdwJUVM0Giil26y+ei3FKDVqjlAKU01E7Y
9aNv0dCaNSCz+OF+PbPzy7Yp+/hPppXpEZNC43zTPaNEEkHfNVbVHhQyokYFYDEEV5V/dWJVWnzj
EHEsTgb5Og0dFatS5DO8iWl/KO+ZT3y870tU80Fq+q+JaVnQlPXY3pX1SLyCCp2WMRVTt/YXejCd
fm/rpqiDGOrHfU4NOgbCssU4fKsd9A5W4Ke2yfyeWTf8ytHeTFTx85PImFK/eY4v1VpSq5J0+Imp
ZbbfT981yCi5G2hzdb8Rh/xzw1pkgmmcBoAE0+g1g7yw6QpCC779azeFSqTzFlZeBOCq/7BH3l2P
OhcoirKYE4zz2zykySB1jD0tan6wgtl4l6SiJCaHY9i1KOAtVLzfsaW/Yg7V/NiGI2Uh23S1cAnp
xMUI3+N1PJorxDS60UAWQBG5rhtovIV8p4I3RhUKSCmIHUoJHxBG5oPLf+YCPaUHyCvio4Hktd7o
anGt0AJ7C8RNkdlwFOpDY0Y/ESpLRrX4T/9w95TfgqQ8kWwCdO6OIp1Vyx7RFglhtnFuBo3fCOYR
xOhbUrfqFKSijWfJTcU8C6RC9amPkLEcXlJgOP8nIjnKhytyT3sj910DRTGLbK3GN6+PqHwiBynt
/BZYSpBe0iF+8ZlULQnuxeL7tAyK9aGp1NHEuCCzRmwHpDJfbfRlKle8rKdlYHW19QL1udzh7ZDL
Ys54TAC7tx7QnryXPwdBRW64jPY7HwY5WcXBDXL7/My+oH1a24DUMszEWxCQQLiZ3Aor4vc1DoPL
nV+mscBTC9DsQ9LeNXIMUYkJ9ojjn7b4V3ZQsqTgCrxvneba/eEupX8l2KjW6MSsHE6PHbf5J6tz
ZD2SCeXTVTC7bc8uCwxAQRb48fZ5vx8cYJXPqJ/sGQlB+mwTLNwpkhwADRooXDo/9mAPW0DLrtCS
LCEJSq15yF7Q1y0vvarNR1WIvpAXO3vwzyntBRzb6F2iopd/88TkJG9Jyfh2lax8JprESA8pqz2R
I2h1H9nGhFxEotMIJ12c/EvdeAYaRomPKmx8GSMYjwNUhxqg+cz1OOGyVYdLErCyWsIt5fR3iYfu
kll0X5bQCAUlrOaxp8nA3kQ6cGA3JCBEza12e+AhJX5Ezcv4vmRkGEVlFPl+wy0Fkt1pyKTIK/U8
Ub0ZRjmPvdObKVB4u0IWwkCu+73kRi/VPTvu9qYBgxqIn887vYYg59jtk+uQsdNJGykAOwSBtrK4
D6T41VW0+0VzBwObPa/xnN+AHvahweuWfjtC38WCB5Pwn4PCjKvUUvb1M6aGIRT/fsApafgckcYO
HtjPWrncpXHS9hkDOwuhJY+2Lj9VitZ/gnIyvjr7G4+qVy/TPYMMGllRfnlu90cedZYToZw76uzW
gpNnJgohSA0d2PA+U3D30JBOWc6qxwj+KNhAryOe0ZMqq85j80qjxpPDA7d0uD2b5sJ88xcdg1IE
LcBRqZa4Tudz1xeMtFUrP0nWNGgAfo9P/h4Y2snp46/nyKgmIlpytsa3PP01UF9PYuKWy+J/y19Z
KhHd5GUOBpFObG6K9SO+Xh6bo7v2QnO8AWjkRG46lpX9y3Br+HgxjWRk6/p/G2S6KHhvpC2rc5Jx
JqimZYn2F5z8RkXCPRSJp7WUIn27oh+y2ZOqfJd+XPdV6zJN/MUaOyT8ooTMx4j8OpoNJCUZMQUB
V5av4Rm34pT6XlPznyeq4Z9ZrEYR8AGF8lyDIRlGDgNV3olT7Nhg/VFKjVB42T5modg2Ytrct4Va
SOGoqlzSOqdbLiLkvcosx13V37dl8g/UEtHQbufSwP4LC577ulzMpAcxwH5HMdetF7H+snoDR8zY
Htj4tPnVQCo/RnXh09sT/op8z61FyvvjOSN6glapW6qjRtzYNXIw7sMSaddnYUAAui5KQ2GHEhZm
3e4rMiRZ6XeXhR7IoXwqEfkgBw9Qja3apeexRIOspvLniI4DrG8FcdJEiCFab8bZptYmEMGgXtek
CSbacIsiJCTPOZQ9tQl0fon1XssjXZht2zhEbj68cMvhAZ0Nq/OPGdvXKfOplXi2aA9k0uOVGwlw
NAePvs6p87TKK8ZJ293/9MWVWltN0KwRcqiwKUN73YmxLYC1gt8r6xTMvWOB8rAgJDTbKSgv9ebj
f8T70SA7rs0a5jdDHaenPdP5vio8YI6ttxEfN1/u5RqbBN50nbGnqpWFQj/J001iNfoA6zUkJrZ7
Y0ExRUBx4jT/88nurxSz3M+XzoRhmlZb4z7j/FP/XlEnG9jAkD5x79wSZaS214O4paki42FTUKBn
ueYCKdCYK9uCA/SCdYScyTCdaLOCpTyB/ivISuvSm+V/3vTWlxQeLkqdJ35mh87o7nwmq2pZjmYD
C7y0QVuPX2ZlXYOOrDYaW7Hty+d9JAiI+9s+H1nFMqCp/4QJMNNrCtvaQgRuZa7k7ixmAfMWQO6h
ltS0Qdhl5FuLgKecfAe1pBSk1Eotxk5+0mGxXqEeZZ6vhlqjdu9aeV0Fc0B5xp7skSdKZ+SFz/dB
Po29PHPl/bBpdNqjPHpVHp82uLNU7+7R7IeG2qkDxg8qjA3s/3dXY6N93F/1ToFwxKf+A1T9D3kc
znl2/YPxPCbkMeWG1d1PksdaUNusr09CjmLQhfc4RQ7uKUt5bWkSeZPPdmQE/8jjFF+XYvc5O/PK
wZp8g4OxGRIe5rLtJa5JRz+8hq81bUPU/uNJuRQaE+l9O3RwuVurcU0idfwP09uI/QJDNYKbl4FW
tY5RBTmhYgtTOzTVlYURHTsflSTTeJ6BNza7Q1AJ6Xw426FOKJ9nsmAWPD7iDz/O0w0VghA10pwy
9pC74hIbZhHC1PRuIjIIA9zA178y66ni5RBsjHK5GU7V5CZCpvnO7PQ7h4msZ3j0kNfWJD/G/JWP
LfXTxkGHGJOYGv7JUe17/kgrBAjvJJqKb+2+M5r8IjQgIFPk113tpFGToHr642SUFZQRLByetIe6
/tEOZaDXuRALoDuvEgDWBbp9gWqcEd5sD9GcvDKoaeWvUIzixnGgj3UenVMIJ+7tJA+qrwUlSxr0
CPGD37Y6D8Q4kSR9OJORSlEUWYDbWCdwAqAoJ9uu80szQoiwbNCfb4BojPI4E9egJW6Lzwvyt7Jf
ihlfEK3aJoqF+GPoK5ReQb1deCOf2d2CAj3hUgTRusYAJsI3vY0XFr7xERHJjQ9d2Tn1AOesAJ26
jbHN20diHjD7eWVDx2GejzJADHd1P/pQk9+r/ySlDoU0pd6MXJMpMBex46asDY08047y+PqR5L0E
rpiyp17d1JBk2ADWKNDHqxte79eYvOlto9jQys1zFUky/OpafMLGsTgn8rJfluePsuqenracX+Uf
toOBJMXbD8ki6xMWzhZUM+E+j2uwYO0P/8S71UX/5qC9mOkn7eJcBg4UrysITN8d54Tn9pTMtWdc
s0WMrxC2/ZoEyHLIrtwOsj5vpngWe4FPm3zNQee2n1JTBvrjo720ooGoCx2PCKDkFPjmF7q8NDY8
Fw7V+Sm14gskZZW8AR/MWUXPcsSedKX8+q4siTtnhWNdS2hmLq2yvaxzBkiIOgh9dNgT/Z+D/JQh
aqjHV3XhblRL5EcJxOKQ8oxOtsUsv4yxPLJUyA5jTyLkq3PiC2p66hSBgaG2Mju9AyuXcGq5XfMp
fp7rELHs7RfcWqNZ+gjtW+TY6Uvf4JMch8TxbAFaYn+GX35nTW//7VBYokJXwPTvPjvGOO/eHXg1
MnQeXnnl42vDuLhKfojsjKB5yXfShD0/JpXs6R3DviOAJXbrgeDG9awj/RnmHsjTRzSO/+mXIF26
yrdylhs5XBI2CR8Ax2ELVsFIcS8iaQhQ0W2oayN1JK2OE9vZWOZCndhgYW8Z+/jYGgpFrQS52Jeg
7rbMCWhATNus63ZHLhtTTdR8cfFNKV9lZNPZwGxfjyZuYpT0Fdf1x2fcHDi2SWm+tT/DwPs9A+qI
7boBnwOq0f6XlbNreHMAWBLg2G4y2zGSrLItEq4lRbry4atXsXh89KUmwBtIB+5PQ5rh4FcAnM7V
voFdGLaCUPhmt2eMBloSnUsAThLyjDvd0QX7cWh/eggUHED51zg+IvARwoakG34ISMRoNehM59lx
qKrcdEDXWajlKpCiOuA28oH3vgnRUlgBHAKWQWvOoeqlcTmYe0fB5oK5bH7hzNxLRumqyWoeGHEy
7W+xLJFl22Mo1AM88c2APMt5iWLwDMg7YbW4O/3+LGWEpqVN0T5rtPOxjwyBJ5Lq3qclYlyiywU/
KHwm2a765kWEYDTbexqEBSg0JCgKtHNSQiNGC1d4bUfROogrksg22rPXjAf9ViiFChKDSx+VuR1C
kQa6Bk2Wz/2grUChka2n7G1UkrHI00x9pV0XAp9ka3bSCxh7Mwoc73vxJ4rF4RmtM+HNqfTBFv69
ExSmcaVpdmCGo5SdOKyxktCEkA2/TfYOfBW9UZ1gKMhU20knLET7iOiemUKQ+qdxIi8lKQJYr2q9
sTLiMHAG6fWeCR0090EfojEB1b5uGWyF3AM3UiDciR5EDjNLiiORMM7miDGVv0ZA1hQQzXRED098
GwBu6oq1YSnZhX+lAlFJDqNstxcXNfLv+NDMS0uVym2CQWS3GvzFqWhJUv89H3iVYpFPabHW6CmI
Ru0lljVpQ/N9y5gkq5go7j3gLIqovvX/tBeU5/0ScLdfq+9mVUhPQM+20A2VXzJE0vRPzA5R60RA
0//0R6aAmNTQCOIS93vg74mJddK4eJJyYBRVm4qmTH54gQtyLjTFkF3O5eZB06hjXigt81CRa35A
PUmUzoHNVPo/f2xpBhbtvMLE8w7idxG9fJeK9q4cxUHmZ28scY1lDHo+Fla1ektDBwKOKfTfPsAt
JtOoyDYs9FiyES5BQ3XnFOaoE5SGylj3GUF1HUbd9wMpv1Lr3Gsvb+26RtV7EmVHrlGlOFnH4Ix5
BpyfYAJhm9Lf21/Khxecqt0Dp7IwRzFRicVUHdmt0nUkthlTyNzXPfaV3omcA7xzdY9YHut6zVD1
VRbS+0VMtoTKq0n3+jA1iAVVE4jF6jghG3TpMZ9f0sDk795LscqaQP4rhzTz65IPyu+Y5l6g2lmh
qX0hx9ictIH+tFULRwzPObjHASI0dGZpdZQR04etkbmdcQBDvf/M8zSMERnKaD8vcWwAXKqUXMOE
CtUCL5bIKQkATiH+h+Vr83k7tMAA8j4rj8a+JBcPo1nuNOXWJQqaAe39+hkRmiXqe2hJg8U1kIkP
SjC+cvqlLWw4zLAUJPe+5Pehj2an482no+Iwq98K4qsTZlAnp8HacJ+YCPfeTpzGmoW2tZdrtwdN
mBjXaemtlrK4ZywyD3vXlkbBn3BqzYiZEw+M63SLNlMhChMBjXH1BxSzINCCNolc5SYSABZ+345T
2rmUu4hDZnXnmiJtBjBT78uH0/V3rSV0BzftbXHfSNrv3svVGM6pzlGRIAKggQlDo8AcRvGsy8aL
t+Dopu4oITzG1PaPMGOrmO+qxUe55ZxcPp45S/5ZoVDfP6ACFBXC5B8RhT45lOmDvt25V8rNZbi6
FqNvW7xe8nyHGJe6ZJiZ0kvmGjXaHs014Ks76l74iiTVEaeJmyNbzDXEtmMJHYE2B6oqeaqLUhnV
2iU9uKxVdZ0ustzvf8vHEDwfIrxozHnjnDJp45+Oep8IYmOy7H/GGgDgcajB5mcU/EgjR+kKkW/I
UCGdqFTyTzRwXczTnaq0qjgN8e08EHlcPWKOIl9B4dw6LORMp9EYJJe/rRDqiWDWM9sUh75aQ7dc
ddkcVG37UwFYoLS5ulkhpXHmFRY7F8U2bpl0auv4f7nP/8ObObKSQ25asFjNft2dFNbUgr2eDJ2f
MYUK3LdpaiXYbj22PjctavwA6g+78hb733ps+5DEzmBS9rtBbd9G9CHza72KQlWPAQ5OzFKNtA8N
T2PIPDxL9RAbBEkSmbk3vniVmfVm8VQhquIwwWKe3Fhp48sOvdEXj7f/5uRdURzo6vFZSyyt5H8s
Uzf50Mr9D+9nlPs+Vhg4ZYq8ia6ELemn1EPrECE7INjxmEPCq5jlPUt4wZ2p/uV5AivtAl+O4hUg
KPKjzcYWN/d5jw1lsUTud6pB8VcSR8ApiYdWPlbiBc1AClz9zjl+0dnqSPtrq6u/tUAdKDwIhFhN
EUStbJDXSJxApu1uAAc6+1axj12GuJTf0EluBNmEd3oCghA9yVl/kiHUUwzLpUlIIgFkpTKbP+yt
aLL8omSLN+M5tLZyXZsMaxVEOSxjNGrthNekKmGWhDtF6yhqS0kN/vwOmfGG9DC/iLMRhUBFLxJT
gubCvxQxJlIXegLoZuzXSD6kuPmUydyFV/7ou20fISGpRPxErUOmt265mp4pw3MdWaOvY3CMV9Jc
lcEHf01dI4lu19yztU1vhl9mI28zWnwxKlBZ9hqZRBCD0qtALp/vnpHcxbsJ0T+Wfk+i32mbS0ic
6AtWWR01hGCj6I97++llMG6eVYTwCOxhEGNI5JRCA/Ydu6Faql7uWMcGdD//M0Pf4unuZHAwrAUJ
ewxpT1L9NmOfgk6IaPA3EH8qZodf37CnlYO7ZKOfvfTjncD5ic17ogFI/jE4A++nZUHng2lruPkI
H8nJaPIT4DM0/Kh2tgyUG4t11e9C69nuU7YUVObRHzFiDQSBtS/+ky7LwgsJw+kbN5CaKz+b7xEe
pVX4kCDxxq4TnzfrwFERERLklEqgS6mu1llkaDs0n6G1RM3OFG9mZ0XS3vsICBvvP+S19msh4UkK
ZQv5TT2EiKOPM6HobnIJyQtSKMzaalHXb0i8NbrtyyYR8tRmUI+Yig4cf2kQUfMGgY675dT7B/5U
fEbx7f/vPVl08g1eZ9m+IaEq8uFOaoDmTvHkp6bUBtOun0xQxBqYcXekJPVJLcXy6D3v0SKyhy0j
iG8oAYXSf1D9qz2gLCHp5dh0b8L+ysMYXT5T88Y7B8wNXfhQmth7GOoTNa6G5wj6lHTGIy5KOBMm
N1jDKfCbzTXI9tXoZuYnA4gWnMKD71r9BKAvrxI+zz9xqY0BWqH7L3y4GIS5ozME3+9uqh9uXPew
/e2jak7ISCQAjI8QRvVbgV+wxLYTpaQEJT7oVHYSv2PO/fIsIYjptHUIPhO1P7mCoIgEHruYX9Bb
iDRBaYMsAUjkt97QxGXcdvy7fcn9WIWpQZZpWjrF7lurXieeLeVMS2nTvOlyDu3PEJKp/2u4rtWp
B0um814HyWS/07ZzOGoKXF3qIcvCg8T0JKRNpyisqhCObnQK4N3oAxMhdp4KpW/X6eDRoCpUpGcO
cKHMSFA2Jvf6n/NF+KjAStPbGZT5Y6qkv89Y3JY9HFSW37pjlC7f4MSD7RNmkcnZEVsI3vIqaD6f
utWSvZgnaaaFMT0yqo/zJrVHsP0ia13MS/KH4qmV2aJNk/yDt0nUCJ/0S9KoD+JEMvMAs0cIpXqW
tmn0vUc4g2zlMuTSNQgEJQqG+/wEnbHL/xrBpJSzETjIBqxiPcKpyXPZrO/1gdwbugkc18t169Ay
cnpW6zLCHMjhYy75/uSojCrSa4faxvZ1UUF0jCoRkUKqQX8tyi14jHOzIL9L6DBxox1gIK8NIy/e
2e7E3X2kusEGc6HiVabhA5g0hQ42phAMZQ1oSZkEyP5fhJJbpQXZKqMQbggcEhs4duWgMGi/0lY9
be8nNuBT1vpL1Pyj8+bq5jqC1hhuyaiwJ9gOcOe4sf2vbAeVSokJKb9nhNic/rzT82Hgd+6/ErtX
Gbb0aMgeuxIEyiDjPuT/xkNMxq7TkPsydR/GD6DCzjigKIrHRypEyamEqv7TKxu/PWEwrOuqtU1z
Pk0LAylEFUnMGfbIKfHDU0dD3Yf1SNhRmGEvzqa2jTxAqEl/jKvtO39LWiHJQWBYKoYjgRM4yVP/
X2CEb//DnGvD9kr4bMrzu1I32jZO4RHrCiw6FNKww7AiCfkUka8Lay68IpGv24KjV0Rk4TH/uxxW
rJQisAFwqUn/NphXEZDJB+OYGKFLlZ7qGTnddGFQgaTilH+S3sYWsYTMolE6qYlIbM8iDuWWyUVK
2eW6JGonpS5B5DcIFoZEJGTbPv33NKJDKFBk+HpPEZup163yRoO93xh2ApYVUCLDoBVWt36X+AnA
sxQq4Ui3UU50VJdORRa2ptA7JSayT7TqKEKef44ySm+805v4V55DSoFG85UyQCcH73i8mrO067YZ
wlBX6qytowWtkOFy7o+E4QWXHu4CWZMi3tIVEv3nUXdrDvFQnRbldcmAIaojHsjisCsEp7UxEMfJ
eieTtq8rwK8pDamtsrmfwScNVQEbbDMvMfw7IQzuEJ3+7SRSVrZadNyMeom7jJQRtkDkr+93/vfh
YZO5eA6fpEExZbc2XMgUQ3IYIi7MYTpNBoABKptdOnhsvScAvcG5d6Wg4IvM3gYnTBj04TY9s1y+
XkiZ3h5TQTXrohQ6LEMVPljcB/JB39s6TFXFDFI+GLhaiGioS4Eg9I2UseuTGwKejrRdePuYJjY4
CfZP05gsHRX5rBWSqpyWI3eE5xC3LzfCqiFUXtCGrk+Ef/aSbI8RnGG1/ag8MiZFqC3A46T4pNB+
b00YapnK2H0hAM9PIkXAvB4Q/wMhxG84euOOFT3CLLidTCyx5ZBzS5xVNZwvZotD2dNMTek1HIiV
Hi9SV+i9UZFndQwEMaNqmsG9js70cX5Rdnma6yE7E/NbHVQJ6VnYy+o+MCac6w+19aN6R45fmuC/
ESF4m2W0FnEOeGkm2pyxqkKASIK0P7/vnTKAR8SbFei2iGYZ4v3FM3/OgWlSn6Y6MgS6zpg+zAW8
CV/jNgVzUQY8OTY0idati9ERrI+BhOJ6R8q8korGWAjcXC36TXBR4H+L/BMf5jYGb5q7a10RVJsu
d4VlNJxmNL7KZbx9E/oTokUV03O7HoJWIn8bFA/b0GQ2uP8skllYHIqTsNx4IfGQYL+mlQellhWW
q0e3w9+7KBhqviUbLihKoQg3OlSb/+zbr9rE+fB+Xy1OI5wknCcgRPnuUoaeOMjVqv58vgDc0qMT
BUgy/GjL1lT0WsnZDLlWhvRzM6gAaBcY0h3hRpV6nkYTjz13J4ftOmQwufnL+kmhxqL50hygvrHR
kXjVh7hmZ+dxPJzpu+UYwse8ioAQQ9HCwzkh3fzICW6sv6SyZvn9z8/TJ1aTH/4fmxSkOOre6rpi
W6EcNbAcL6RLoyFyFLHxD2eYpNjpb7d8Ujb6snqHvXOKjRkRS7IGXo7ijH7VvxJWahVP9IMWgqzh
eKpgs2brvil2dnpr7CfW4NzUtNCp0EftXUAGIsmuKTWcjrLvqMcml01XGn0+DqI08Q+h3lfNl2F2
ZFsCCtAFf275QzP8Q3tLWyEPTDF/1DF5dG98WzQHD2qKU95QqklWj6wpdCvytuHTH4AM7sl5GLRD
TkKqHQAmlOewiF0QSy09jLLtK2L5PhZc0GAPFa1PYato0aXI5o/hS8i9m5Xujn9yoakR56qsXtCl
i1mf6t770XEbHxYe589E8mkAEOdB9Z//6RK4A2kiU3/mMSKiFisw45UnQKcj89mRy78vZisTrKp2
E91nmaTTAiGo40p6DUPS897rffJnIDZBVLgRwfp2Wj/CZdlOTIAuycK958JzSGUyqeAHQkmZ43vX
XAfPXNDsUPwLwj40sfKqnZrkK0/IOEpPjDhtwOwes45YOqZqTSicw5C1fQWc4yXOT2Ko43pjY3XV
PttupMI9+flnilDZfitkKuQ4COvIfYXm2GWX5ZW1V4HcadwDqdcPq77YT2glB6oS6wxWGT0I93M1
4kvrwOJSijkHIZgAUhPWdjQYPghlyROmVhIqR2jNUc7a7OqUDwEtqFVsTdrbMP8mw0dNA5Gtaiz4
tGtEJndw5wDilVikvcVZKGApGCS8Tz7UYsowCrvUKHSRkAzHOWYz+Z1V5C9gwKVQUqRzlWjoAroJ
f3o+645910HN8OdDxNlnvQ3oVQ0xQxR1WRH/b2lR8cqNPdkptNbnDz4+x17Tl6LW5GFWTLqETmAy
XBFPdmEfxLj+WHW0Te8RdJl1mtLfy7gZWBbMFPimZcmUaVGnNRukOvqqq/adsHMxM/3aJjc5WgvF
Q13k0JOeusx0XdZwktjD3HRn5V+nOdxUh8oN+ARVF0vHs683jKjOFVlf9YP/DRmY6j2YTydU2WxL
8LPXiMahtRAUhV9ULgJ4ffdt4gRg+WR5MQYuv8jLP+JP8+znA5WXitVRBaYHWa/cpj3qEw4/daB2
Erp1ctlJ14eMk2ks3SJ2fbuM9dnOki0SE3f8tJNOL+/sRhBg4YE1FYkFjrnD2odySk9liVLejUzU
kNDZS0W+Gt+o8/gT9doOqCv7cVL3F5RQK9MXHVu6lJyQZZCGSNbPvFw2B5A3RuTpxoGxV/gaQ4vW
J9qt/vwk+DyzIbeNBo5dXBZI5k/ASWhG/H2X0+0rGfgzLu0D1UKnWun0iOYMUZtjsU3sOTN/dX/G
fygnDLJ3L0bR8p42c+nWQz8iHHBhxZqm+sUuRI0UOPcOlzIYQuP48xHR7BN44VfP681hL13tTSan
sVWsv8RPSotwBkjA3Ngr7EtAkZy7HcLWL9l67FFKnwtc5oGqb50fOMdvcPVoSUJVzab7E0n7Ls6F
q5IOWttlBrB3fIdCU7chH5SyhXwicsyCFCna3td0VqFTyB0fsObMgIAJTZ1JyGGRSOtZeFZZlX5C
MSnj4e2kd60LXqKPPVjDB0Eqe3dbnbBPUYgOCJdkU7ggke0iiq0SpJZKwydW83eWzXkdP8prpqHV
ZXLkzpSK+cMKov4voxHP7HSPfO4wLL7MkxNF6F2sz6cKuyX/XBP5hOaOns2tbg5ZtLReFGulFW+1
lOAlFTM6LxdHCavXlE2zSJj+El6QZcMWm9C0UWyTGn6yASguwMUvTmvXJOyr5aDtIURgfQjUxTJ9
4e/VgJ8ce3sI2/h6+GHECo8zkHkMBhF5yCK7PweugLW50LZBE5EDyaJ4MsRKPvtzfxlyC43LfAtY
JE2EyUjkoaApwcZNf9QE0qV16OQ9C2iUvmSQB5rqQk3x9YT41l4uoYos/FfpQTwTY7/QOMzjI+N8
r4frsPS34b4qu3Y/YIcQHZ1XTCFJDU+KUtRSkDkk4P84OSr3AntMCCxPxKamymeoAt6JXHP2Ifwz
4Ieni28DWk5JdmMWL+7Ofs7PWX8g0EcvDrlPszV7ySMVmqpVOxppdzMCJvv0F9mTJHOu/f4kEzmG
hc5w5pkbGkiK090jC+WO/OX0bfu9mLAgjpgGwlFQfhc6htG+YX9vUyUb1s8Tae/PhUa/PwSW1L0g
RHBidNjXE3EkqJTBggmYLSQP7ADaRXomLd8q+De59UCwUKqsQPo3DlglgRnFXMYzbyYdRBLtDRSi
3cm8zWBqwB5L+/H5WAuA6Tu/9NqltYvRyKZfsfL11/gaAAkAavpMAoq/okvyY+sWXgxpQW9FlR0n
8L6wkd5jnt+EQDv3WUWd6IhML/uEN2PtSmlpDq+She5qs899mQHXAsHI6spvAw/F8d7sUYgZRlzt
tOUmHbFS1Z2/qEXBx2/hferVB7wQbQaOFQ2ogc5lDNFCaz5EpvI0wgiC9+RVIhfCZp70u9QwGFxI
ANkha0hu+lVpKEGOiDZdvUH6RDEgyfGPmqfL60yR/XGgPVb/4vlH3eTi18KQ9odmuivCC9CchmdB
FaZy8XMefBOp5qnAZaAvF7UiHNRsgdftpNVjEabtKC7fp1hjf9OrSmrmX+DLz8nfC/um6Cp8O8Zd
zyeAGQbKm8ii59U/i8y5wZZEPF2dvW3kIPFitI3bHC9/c7mt6zEkFH35We2ZbI7ZDA4OrPPigwmP
H5l9BA2EcXwRsgWcoV8DLeNFqY+XwCzKiA1fQf9lnr8eIc+GFv2a4v93mE68fYy6PEA7WSaLxeko
aQq/ONhOX4LUekcaCmrzN5rNwuXbkBAeoQuAid+7MY0ls5uLNdmJ6EkziiPji3GCVa9AuWWUWkJL
Tnzq9g91D1LPvI63T6H14YqDuyZP+8acGb4N2p1q+JHCHE0GdFFCXgGkvk7oJyeVyY+oVVWohyYP
IXrjGqlScPORVZ01hVU+/KsZAIAzMJdvaqSNHN+1Lu3QPrs5ycwu9UXyMAryeFH3eXPh1MOUfRGv
p9YJmJcC01i2H4odt588pj17JLlX8DhyewX2BcxFyoMyIXAwxNxVypAm8V5+Oct9WRKf53669nkr
LZlAn5iZCPnhVga5eavwpooZLiZ/U2WdhdLkmOp5qK3Q4z/oCcac63C63AnN7HjxAPBtEhCKKeZU
oPeZFdRqVFeSf/628A7MMr+NgmeidUiC3sJmf/8szd0PUqfZ5Ae6X0kLv2N6laVgd6EEgbK4Wpc9
COE851b5UexsBHFzSlRHZec7JSS6LdrccW6lyPzjzD5TUQYOjohX6qmUd7AdQWR/eL96rKrUxoe6
/t2IHcaRQje0X0lfp1XyYEHLk0XDMHqlANdi2m9XiEZDiFp6k+8dVJ2/JlROo2qdPZP2uMq6Rr8J
OHYcO4k4atbTYHQYGfWiT+pxNY7DupGM/kwL7Vr72eopDPTl+IsAcau6UR0h17fGwEaZgFeWmYZ7
y/s4HHjEqJkZlNuCu/XmFykhQhU9uHGK/90vWSrNAo3cZDp3zdZ5FAjwr7BXakNcjKT+l1nMuxc2
f75/af1lGjZM4GsXkzAE/vdx9XF+HZ7HeqpbwJAGn564GdYRlwQBgTIg9KHaDliV6ffWYe1kFevS
0SeVpqSY73QGu2nmd3SWvAfvP1MknjC1qP7HyXia2k8I/OZiY31QMDq/ItxIqcCic0VuTY2936M8
xdqKvJrXj7Qu+2p9/vA7f0v7FaIa7K9qnQKFDNKzWf5Hjavvt5ecWFGUa9rYLUfz7To12xKRkoUN
cRWSvoga+sg/Qd9cX1yYvSpEepccW4YTRlWoI4/zMuIqMmZvWMcM5PzG5rGfGdJPKs1U2/zgC8Gi
bd1OkCZ/QKT23g0/FxjUsV56TPOxfm0JBAVh7B9oOSjjLLVv+Q21hr9SfhhJIGjpdIzvIhIYs/fi
oduQNSnu8tOi0Id8UWD2KiDHxQAIvGb7aaJisP5RMuuewXM6u7s0Bn3bFVhWA8d9wFiu3c0npf/i
IS7ozc6EZe8IijBgakpzRxARCJhf4wgMZd9aUysPL/Thd0vJAlXWzaADFsAmOrNjuOgyz6mmJc1q
5MnREEowg9KIxdOkA1MZQ7e81mz1sXn6XrIxnh1u2a35uivoEP4Rk5a16dQWG0JEfeLWrB51Lr3s
cNnJlc4yUY94G08FoGk1m8r1gOpXXJ8LVa55uxdhiGJEdK7cI1Ih9EvknwYzd96qpv6C4O/1+/3N
Uk6Eu1dIZQcafQORmuVWcGoWq/TsSoCYailN3OP8aZCoYDspXYSTtc0/EhgYTyKQVM0eiHKwh0y6
65SJ+FOrBZ7WGGg2kxakB0ZdpFoswHaG25yl4vq6wnEUmJEx4a7TLQLVvMRPJx9txmn7yDTmPdCN
fK9vVFk6Ar5e12JtUtCW4tvqUCGkEcyzYtGa74QPpyCwl5SjMyoJLmnho+7ejlbmfU9lgGP6VbgY
KYCd4Mf8WiJW34A0bBoyRfTpch0bJgmXsR4PJYFXuvnmvgPDsxw1EXi+nYMs/NvR3sCSpbBdtvtv
F3zmEjfZcKdynYXFQJrgxK+wF0jVZFqQwXC94sQfDYCjpxZG0UP23pgklfx12QUITuA5H13Ru9FC
6CQxX2jz+1OvphLFtyRDB7WI/NJqDQS79GxnqaP+JZqq82ylgJgGMY/yA4Js60UtgduTmEV8gQOU
DwJlGe9zFXcysHeLXWHDt3Tztc3p3nuq1ImmPDhXBiKWx3JF1BXJ5Ffh+QdYv7DeNImeeBymaEqo
o6aV3KqCbdZ3sUaU1JkLFyXz7Oi4fi9fxPir/8d/16wUtNJLSmo968rztskcmBdDlg5p4rtTLLXb
Jw9/Ja7L4uMt55AgXWf3f7hxS7NKpylRUAzQTKpF6urw94D5stU9L4GdD9UEvV2ad4IgiXXhzfZc
InVwz6NMOb8YHvG/DYQGdNS9cItD1w5mz9NhveTOOrtuFJOL7CdTaMiSaHFfSDzQFj4Qtyfhr6uF
WloLj/HMVeU3egtj5o8dumD4aj3xfZE1FsQsvoky1qSefZuNe3DLEmfefIZqxWBE+Kzm5JmTAkuE
ZsmJPenF6efMQPocbx9NmNIcnQPVP5z3o5dCedeu9y14jzcpjWBO3BxGk3aFRxedFuoC/lqRiTJQ
WiNeEMt1qfCwvRm8Una101Temw3z3q2aI/rPtARoMDMwXARK9nc9+HDb2hWoxvrZLD580DYJbi80
S4DPXafM2lJV6HwyBEt6izrUCxlLCBjnVSXl1Kc9ld7IrGIlNyCT25/mZrKzKSXCe994bbkF8Bb7
3Jt6jzyf4bt8Yy/fqkJDFl+IIHEBY6G2ksL8b9CzEDib8AHAII9Y6p2WC/em4yq/IYunXLPHC+3m
7PwLbw0L8FVgF09JM2y5C7Iop/jxW9XjzU3sNfKK7jVr0rVDmVJK9WANIeuXmIi/HkuxDIREeTl1
RNQ4NJVoM0k5T06xeu+7O3PNYzNV8wQQ7EOk3x5dlv7a6NArqayrhax2zIrmHdVNd1NUeHn2n3P1
1QAExTV0CcXuOAy28/moKVhSNJ8eGsrPwjoFLI59wz8YSZa8YoDQ5WNjSct+C/XtQz1QKZnaAHSf
dHNU7e91vSD5xaZ/GnWdd08YFtO8cGpJ0yNjU0H+PJlkHdj8s/H7hw7iDTlLsH9bXpd8HzQWNcwV
phaXjBJqFPZ2pl7g9su3aFVeBgv746kikqDgI+UeEqv8BtfglNfuwRoLf1GODoMuMsBQPDcmwMzs
eJThj8v4mOg7gE+wtlH/yuHBX3f+VfN5gBLY1ZW18J9hx7ZkmeqOraWl+bzFi+KjBp1BmIwxsJte
r6aVLOHutdaVi+NETkB1NGlfaH0yNtkpsnt/DS56z4FHWAdoTFK5A6e6oMsf/IoJ4S7MevAMxPCw
KFtwXk+le8R8G15rrMrH3aB8xroUJH81q1gCs8VeS1Bbw54pHfDXjzkojawWAZyUvCNdiFVajDue
qyQ0ONejRs9WXoKatfkrdZ/0afpUczxuYtzcrbv2KsiMv07ThuIQbjGPc/Cf/vt9FgiA9UpB34gT
sIT5Fx2blPJPXdQCLXFJ3Y/CUkoclEZXmjkB5L9JCnwPbNyqGoR6uO757rmJvUB5KbUDi7Ni0pU7
fNT/oPO3yD0Tia//nKeblHU6I5tO6w3lMK8vMCuwuHgZ7KeiM36NnthBpBP5gQ+KbxbSrw27HdS+
nazWlIOR6LgLomIZJ7H3Bgq6PADE6a7hbQcd/mOtHTMm28mLjnZxMVkiyijLTwa96uF2VjsxTXzs
U0jV4BI/L9WOEKHEbczbw8K2i/nge3mPVAMUGs1Ia3HNbBIQyTUDjtJIebbk6pIa2L8skCkuPWp+
+K1qSPmiA6SjPG8ZJL4tC7baop5AaTcbCVeHHftXhRUUNkxzMFdHElx/9bh51asfQezz2A8TZO33
m6sDweJTxL3jo3QvV9XojPzDQYpA50xOBT8ZsMDWQY6gApKaH60REONwh9c4is6L5cleWXYvqhY8
i2sTzC0fNuQj6w/CSOUMCwAJiDEhqF1PlDuG5z5w0Non4Gpo1EkJ1UtCeG7+f0RLBHwgimNylhm2
otJQd5VDCEj9NHMHuSR3idAD0AFkVkB7aMgSOoXLI9D4xWNOco+O/V/K1M96CwBHGW06NG4wvFLy
Ma05M16zU87qyetFgFj83ZTtO1Op4I55ggw6YnYXLXEhs9LG/ldyNjZ2t3Q7Bt2RcE3xtRA8VAE7
zL0/JJtJWWhCdCoI95YUFBujM2npI2U8Ufe6O0pmobPaXTxAOjNHPNPhXOfic6p27i3rBl79GmaH
UwAltBqVGQJhqE3HR63ujXq3QaViMymZtXhSq1uPJwW/yKoA3eK8WSgy/JdvAlB0p/syfrgV4O0s
HCGp/ogtdpFeOo6wsr0bWNexTBsOq8yPMdwaS2xATntYvHcqZk24FYjGCdhBj8L7Ah1lu/mmExHT
Zk8uyrTiy7xlAoSe02Apzy9GE512sIehT2shZsPGZeeMHyUVp7PLkT7t/qDUwDX7VE+2V2hr9qER
CpC91WN8epsfFFymTn9NBkTkT1SBZHmhE8Ng13GTGRV2FBI4QWDHjJ22xJ/6uuffjiAB3sTrNIem
W7OXZW8H402ZdeO+aSka03EQE9LJ+MBnbKJgkN01z0AaY2WnSJhQyKZRdKLohQ0asp2pLu3fk6Qc
ILA61Xijz6MGfW+aiYLYeI0EK4rywafeaFxneBn6Ng5GnLdFXHoCOw/GEmI9MC7EI4Gb/VpC2Jfo
0qgpiWwTjmiWT24pQQrak/POxw5K2uzEV74ELSsOb7By8hkaMcXV1Zvp+S8cKi0gD6r9KMl6YhcE
dBT7Y2NvsPbX//18KqMQj/xDOc9XwozCLzp2OKRn8TR9cgUKQ/xj2/pz/T0SMqoDBs9FYAJUHntW
xkYms0y90IvGtaL0C4K0dpxjVU1zjaOSB/PGYHnnxqeRRVvaX0ZLNCrOXi5yDuMR9d3xcU9t5K0E
Fn8Z2ClEJMvQiyoAYJr4nCfNT3d54JavBAXSdZbfyluTGfZ9sijIbtjUwsJqVDnRFEpkOFd5Y93+
ZwpxrykOsDA79FQZ33v33VHppVM7E0hQd9smyiBSOHchGM8UJwJrgQAqXh1R6Vh6i3SJD6r4+CX3
jyCWpcg2eu1X+WyuwhR794g4tH8NUvIpJSJPmIMF8z9Q5EwspeFxwqdYmMGaGzTQEVmSEh8sM6Pu
XsZHYOtshyGFkjQ/Ixi3SvdF746ML5zP8kHRgIwDj4Fuwlz9K/YDna15QTqzUi3zRNtlC0KTK+LI
RQsbX266bcU4dDGdSIItUidg5p+0lbwOApSGD5Cy0bScPK0UVI1xMeN+HKhJO96qwwrLXi8/rdfn
avyES380bZ4qPM/cySe/pU66WTSlmj7oa+MJYLBW1FLmUtBmFZ4pmOT2la7SLSgFqS4irhEeoo5H
Osrz9u34P/+F1SKYmHoIVgv+43IwX/cNh6uydHJ44tDWPrqmjK+4ovCSZaBunqgPtJRx6Yzgx3am
Ph3Xm5J8X0+fSmcVeHs4Ec6hCpWy+E4DrzG9RfBOl5xe/hGDXrMiZKx5u8ZGje+Equ13shJJd7mM
/Csrr2/2aYT5WElZyBYtzlOUPJOKMhZgLyAIgm4bgtThLH+zMUqn/wAyVDepaiMA8zENRQWuVdiK
IJ1g0cKrSl1GR3iKR40BVXpOQeEuMJ6sx9IAIKzre7i4Bp0jognE/7sFSVx5VVcbIUb/ONz6LAy5
aT78kmGZ7OeO9ZFEqLP6YGHe4ogDMLodaRDlUCsek0O082p4beEg9OHyjlZmba5Ww3cKHjf9fE7K
WN3VLh8Waj8Vsua+I2p5G1/sP4Cq0bvkLHj1DqSy9DfvPhPdL5l5Z/vM+CHl0C+iOizuYC04io7S
+7uJfbnmaMUB76Y0a458ZXMCmQm+S58uTDuiuekro3fifkqY/nXQfX5BEu8J34Y1rTNpeGrF0xqF
nRFexqSM82CkZ/09/4zbF0ZyBb71nMHIwx+rqZ4y+GFVZhPFjYvFHibnTYF17FjnIfppaGdx6MBw
ux8vUi7NJMq5Rr6jmxUWY2EShCrNzIvOFlKBNvXC74J/LaOHs5sZ5Az37rbGCvxwPeaOZvzsNZ5f
61N6yZ7Mks/MLP7CrmjQUD+Ch88aIKcdqjk2t0h0oJo9QIHK4MmxnZtWvxe2d+o4SwyY2VQhh537
fxKVE1ydZMK3uLwpULgKEpP2mRDNdrDD4D5AbW+KFrVJgAgtlgg8e3VPIU6F/nHXj+mHPWpaq8rx
x9oGc5d1LMepZsVmeCeN6k4TpdJkjW324lymUrpSg3YkpIBHHDJtAEM7roYPg0NHrQPnEteVXkBo
qp8hXyztfVPpXANvTjjv/rt/m/Ha2apr69w1aeoSUAr3mICR3HeTtC2szWGW95QSf2aHLRLCCjUG
my0c8w0d5CPLK3+ARGrx6TPJcvjd/XrmbeFgu26ZlKOuof6EdeAATzmiUpzpImkbkbvMo5t+umeU
G57tFlLRCZaIHwITHqzFbc2mdSI+JNzJ/XrO8kR27/dmKAU11dU+Whq1/MTimrE5NAofGri5YrnQ
ZPNb9X366NhsLv5z9y/UOp/SVJOLzvX0F+VUAzfVpzzB0H26XyRqjpb4kDRSmJMeUlaKITKTdhX6
zusvMowoL04DJTKpTO1/QEzntS5EH+kGPkb4bHFyoorUYTbKb+ivfCAmph6y+SEPk5TSSsLJHHpM
/R/WGkpQrMRdqaceRBLB42IowQatj4e20YJIylxoA1B/4ask1Hrx9jq2rZr1XmXHNOWwFyskfhac
YVpm5RH1Hy7YBNqghGGyD0+ceFKphWb8F9zHL1iBVtPEK9Yz0Po6QXcgXjknBBbTlV+j4fDO54J+
Whwy97i4yj5E0epvIPRGtGEhB8raWVUHX+uz98mWbbVJ1OdkbdLizGGqwyqg1bqgKMB1f3k62hJO
OXv8LYUY5jEJLRasbvB6mYs83Ey8NAZHjWAMlqzz0azTdo5Aq90+9w/GUPetrGUV9dqleYMYbaoe
9PRsR31u2zAoxm5panRg8c0kIRV3ZFV2GQh+CjeTi4NBecDXHIU95UiGdrSqy7DlC2NRAQb54SoK
qx0aOMzPmwp6AMElgYHcKpYXCevLHq2fNZ0rZgI3N3unsJIX0b/OKFz9Ik20qVH9nrEDSTvQSvv5
h6inwWo27tKXPmgLXoN69k2TI3VX2ywuYYf2H05ukiOF0ny6ouD9RkEFwizEtocfUr2ZSqYoVCDh
nmEKx3qskmlbPUzA8liiI5RajBPcoEX82lw29ZLGSNzv7Stl7irpGaqKmK9zl05I4XIlOfcsPLSE
eLTWDGeJFoHQmU/rlOI/DwMmN+SqNHFv2ZDgcknNxdk1+iX31zodJz8lmcKmb1L1ndK6L/AqaABX
P417O1j3MU77GbTxEalJu4SoLTL4b4HZsnMp347rW4uo15oi6XjZUFk1Qy3Tp7ziWbTZQU7SopTW
2CI4tHB89ZPpRah1aKlXCFFYWNnoW9XCoV4KcfCMm/2LeX2MHk2PTzIJPoiJEReY5Ej5iCdGQQvD
cSWvBLFcNg/cxg0CdjC9rAcMp0a2ccna+ALF7lln/HAA2V7CsVrc1KRhYYsun+8Xrs1twVFomZjb
h1CGMB6EOPvrRAHTeXboD/M1Ld8LHN8ppJfai4O0SVqoer7ih8PpyY3llOuS6nUOzSOedEjnjT6z
b1pCFwr1PinzpNhzyu2E+KuCArsxslWsU1UdGBLB/TQdar1TP+0ymEZ0jz00d54b47OPyrH05gVM
+EZXdqUOV6nQq/ny2fDz14kk8ZnvhUgepEMYu+BVDF9FWzgn3V3BMweWWNhPyUfJKz0wL2spO/uu
PteqdCq5fUyF/IY1M88Cxpvm3xL122xj9TNIhnyda0URZxj0iTn8gl7Oc+BApZTnSwszprBnvblh
IPwc/4ciPfw2wQy4gh3/1HAp6NJOERnYbiQopIKIeHmn9AExMuQHZZXCEK7gvUYW3mVKE2yb+APG
xErqP6qbYRdk89u8LC1U7v1E4crVWpd680A1x4dFnvvSs4CULroCQPOip5iFeYsy5VZlRLmLwW9Y
o56I7yDKS4Jih4uTvWc13CUgiDtiz9cC7NhQDWcxep0VOPBp9WQ+QoxMbF1xfOHhcBlonxrgp54a
5Nyd/40yMVYRxh4rSSGkYlXyDDwbViJwBKC/Icef+eMCoUmhZM7vWp104KAbUbbKvYtmPVJJ0PZ6
y7XEZNRiDFn4SkebylukAHISedNp/bn+eE0vB28/+PPe0OGYcvXohPx1FNkWtd4CPlvmecAmu0Cw
qd5oSdo59/CDv4egkPvqHXrqalgt5YKOsasTfjKKtAqOlIc75LW/OWBkC1RGH+r5fLZpfrgTYbD2
qqykdoo/JZATk+pX5EY4sCe3fCj9gITkKUJdh6mGrES6fHmcLvvqQYrNTLVrFCWwhy+7fubZqnz+
noUC6l3Ox2MiRNrij1dJWWI6CnjXErTbKbkWVd/nsSNeTEvH9P5/65BqwfrGU6awcmNXAzYdeLjk
KpCi+Ub7v3V9WBAvb79m9y4LELh1UdA1183YLS3M/88orUiaBtRyR15zaNxRasBG/DILWkiygGsx
m7LKNAypd/7VcJ5zN6XbCQW1lIju8SxaoRmrtkIgC/MFzTRplHsdJVVOmiKIGKDcJTFJ8D84dUPS
g2eIu8zKzGsPX7QnU1LsZktsZbqcl1/0vZ/dLnmn4KBFPqvyarQskSgWvkTKM4wRaS4efhRuSOI2
KmYHcvxfEEzZgJmWPkFcxUMY5zzy9iB6bXTY/9Ddbd65m3y+ZZMQ6uKCe6pVVuCHDlsxwYSPEjuU
VztArx1JZ3Gw0tToP7N/qNpJlmRyZViabJFmw9ROy40efKjw2/oOGHmY8LaQsEY9e9kb05yelnoT
Dwjw77eBaC+yb6mbhCynXQYB9T+3Tk3n1pIYPwoUS89HXHIMvDGOBZTmvw2RWNFh2P+DHw0jUOJR
lcXgFeNF3RCw4efxgpqjSGYKH63w+xbdPqKXPgrzVBPz0J2X76geTwQ9oDKVe58Qvny7ypqLmPmQ
nBfNB7CaKtNEke6uOUMJ2i71KxaRuSSBwfCn1WsUAn4dNd37tZ74nHnCUy4FIAfmny6RjIgv8ZTn
AP4+HkTqe+Dyw3NynFf9YYdfch8xLRvBtS8IPdn7JqKZQNeCCTe7kzCv9h+K9hYEiiywoJGLF52x
QbQc8DJVk4+qDenehyw024KgHNpnOC6yg5IS/yq6BSoyW19L7EkA38KsuftxY3NfDYSeI1cU9i5+
PPfPwbwI0K2fInnzzz0AXQEWyphnbd+cInx1ozEKqX10rnoVYjA6D3+KG0aybDFqx1hugnCFiP4Q
c3bDUOLiLJwdHSy9EE8JFZRNPa1PVddjA0CgNh+Y9c7N4dnEO9SioQwucCx4nEZRCueNL8VvqmvU
4wUNA5vEF8/jy7s+1D6jUDStrJE9qAwj3sG8cBvqFN/0p92NJDGr8H1K5ozcGvwWViNi/BrMiiTp
kuTTWRh/2x5JrW+cwOYje7J6+3iStH3Dig+Zxr968nb0sjyoGZFJ6PWVApJsF5R/uJWsMe6QsyCW
Gx5wR1QtzqFP4MffQFew2Uf+g7Yl66z3yGJdStRYdg7sQTM8dNQsC8iwCZrS6YTTNE3nop3LnyLh
wa7nyErjMlPXY5SMDQsmGq4m5mARuOiYMvLCZlINyIoSHsjPPrdb0p8bO/kPY6TohqBv6h4CHLoz
YMjhOmQL2bK8Q+QMiZQXyw7BjzZ1h3Yt4szxHuYmEwAisPCr660rxeMcJ73ys0mw/O+nFuiUIeJc
HWsOgXjzTVyMAqJcuzddkRbwZd2dlhcLxaC5l3WxVhSOPiTtiTkKQOL39IczGKZXG87R09NS9hj0
IvuT22to10ypzl/0s5uAnMqrpfJ3m/nxAe1GB0eCisv/oVvVkd5p6vXXNHqJ8U6EJBTCKV4B99Fb
PSL9nF14dfAtxCaoZXr7XEJ7n5GYjz7FYk2QhAc1qLZnSSa+G7BHJ34t9hEYrT/iW/aNZ+rCrYgC
YYL7pyzX7G5U3eYK7UnVeCD67fzmijra4SJtXdjfKGv7G44Xy4J5estba3YokXF87YpsFcp6P+Am
A324okAbfToc4b8xQltKWWfRaQTNX24j2kkpq9eUT6ERsmhlM/M1kYF2o5x2sP78VeOcA7KzAdu7
43ZviZgldg5tErHeRy64wdGZ3ajPAHo3LWqXWlULgISJ0Fjlt7udkz4EhYoYxD+O4rTS2AXtGhHM
Wj/EllO/hu2yM88jJaRbTHHBCz/HgsUE7Du574k4Ak3wLisHJTUm6JZF7nNkaAu6FZfMgAnF2kMs
+5+WYE1fyHR9MqE8wxwBKaqBXqhbns6EUJgsxaJfd5WnjnzbTxe4RJYS0nNxdZ6r1EDk3CKVmnIv
002CaDvk/P8/RjVkp1LWchSE8KsRfBCbuEfQy9uzHmwm7CsswfzkJyLjuI5p+1mBiqDHqkKHW/mC
hQgvdU2zPIT+/S6pNB7k6L/US5r8yEK8gBs43X5j/GQSZQozZNrVX24SiTV8ZIR2pdAIzjTMrczI
YwCwslA39qlBHNDC6GS7sP2crhw3Ud9ULv/DArG7fX9SKLq0Xz3b+wap+OXArsEZNk6oI85tfgkz
pFdNSVnFmm4zU+AALrmNS5qCCKIATnxtSoWI/+sdY242hcWE2ifIgMJ9+PzCPbhJ7EgV762CeGTu
qM2r5U6DZxtiEvlC1sY7bqHccLgnVZHAP3LpLDSYvb6V4A2vQkbU+6Sj3G/S5jCRmArM3loakDKd
LVMzkPJGV8rhwqQT/dLUtPCwrn9Aj9EBBaa77iZ52qy7AHsg3KXQDt+YclIHg1Ct5YCk+MAVnrve
mAGhbnUkybD9nMSY9gy3vo6S+XDIl/ddJmhWce63TPnHbEJUo0mZP46nOxJuoS27PDHfqU8o8vw3
6SFRGJwrf5QZtqxTsQgn54l2exB7Dpy+AiqlmGiZbmXsbXtY/mC4R9BJcg2OgDwoniVWQX2tsdiw
IuOuRHQcW+eE+DErOw84rwVUGiGO5fq+lOIdQ0J66I5M4B+mWy6opRvS1ZueKiY80IMGCZ/N6k+3
FSBoCffGm6xFFp4SrQgFmRqFtXkBSvrVErs+fkAI+dOnn0VhaQ/Ump+Gw1+NHp2Z21WdNqm2Cy8l
FMO2o+MGAqusRks08PvkoIiCp913ySsW9LXFSKFx93xTFykjgbgvxyiKQ5JI6yintVsHloM+o5DM
pOwTdLJbG9sWISLZ4kvU5cmqciSYuXjTwPbYl8Yu9AmS7f1DvkZSeaEEwFAsmxeBcpkRcFpyK0Uo
9ILv0PEujhRlPa0vpDZu5Rj+SX+1BP5dcm0aFXxNW2e1nO9mimxvrUSlbkaLQM6rqX7nSAkIeq4X
2voxQIG6QfZozJU61fXAmLVP36kOCITSuV4r6w4tBZxir2hC44kmVAHEhypT6kKD1pAFjdZVwZ/v
T9Myc3i6cb1ERTEkyLf82y73RSbcYtgyvrZ80SjbqgFG7Je1SIvQyvJFcbu/zQrvtrn+x3epeF3O
VkTjY9ttDMv6dlW1Y00b32vyB6yGoTUXb9OMU8RMuDaGCB+ALxc3hx3ztFFtvN5W0S7K5S2ED9Ck
ghktYL53z29qkLZVbztMN83csTaFJrRFyfcKK/5i0rLc+/fYrjKOks3/9GUJcrvu+qlDuhfZRjdE
C9nj4aF7GXgqRNhX0wCyb0eujMaQjxyxlSZVbS6ELxRjHohhOdH19ic4SoV2cRXBsdm1C1mSOG8O
b395lGNAWd55YnKYIWRuLodn5YbSip1XqHc7F6iHIZ5Vacv72Og3+P1+0Es0YmnHJ+/3xBrP8Y49
hiWV7SN2mvBZdqe7hjNNXuj2egFX2jJrz4u2JvWRjUglcuYUkVjlAOG8kRJSCLWeVC+Ov5m9CLqu
76zNnDm59BUBJl6oOxVKhnyN56ROraBTRT46gHBsa345RlmomwCQ5qreQR4MhO46OnrxoeHk+K6j
A2BAJqHlHLYnMIWfDv2KV0Np8PDXIm8L6iJagEJjfyPVlyDAxNz6DcqBWmm+/yc6W2dW6E4tU9hR
nKAqYpnQa5GCPaQzoN7gKRJMk6lDitiYgAPWxje+BqYeWBEjeAMfbfoGRZ9eVU0prGGfwhwtAoMS
wcBDkTQBHLjSlqvZqYGw5yDFuomuq0N++28SCty8ukPHldYOdgFrX0Aj1tciVzNuGm/BlpNpzlSb
RRSbzgYShijzmGQiTpuiGp5bEJObuBsw5owYLir/burA2mpzCzSksvMYJO7ZMAcYujtvjcPgiQOS
eITFiOywusJM/TEOo9RqSOvM3qKdRTcaVPendRFuo+v1hCK8E5p+HYFPOecbeJh1TgSaaakcFi5p
IGxY0j/BVW25xZCEmJg/dlssqcL+tWg6sUFEMM7gtM/B9HtsTeXN+cv/3JvACI4AL6j8DVf1pj3D
h7yIEsRq9QjXUiwtwlEOWqQXnmwTBa8PwW5C15FM44Mm1Bpqzvoky9RKvoYNXzJhefyA6lnkCX9A
Qs58Bt2DMJDmWdvRKNhoeOS0tayaP6k9lCdFgP6C5J35Yla7fQlCwmXeUdrPgZ7Ux52sTPpchb+2
vQNWUC/9DhSI9/R7fsKdoSf+CLdLIDfJWPiA6G9Upp2gKm28KnLMg+9coU7hylNwhv1ClXkJ0tmi
zjOMEkhBupLQ0BdXEVmvvjCyPjDhuX7YiYpdlOrfcBtTeniG429xCIQPZIZs+JqT13l6Tl98Eeml
PqTEuZgG0Gm0eUBy1d2poWyflEmgZadna/xi/CIxSRBgvMZeVMI5rZYb0mhvW5wYS1C+B6zSwr9k
pjHaU06mjWx4Hm/6TkKFNpYAZI0/wNZ1dTESFLHtXCZm22Bb+tjiuyHP7VRl0IA9RU5J7VNMEoGK
0iKlLn8Lo+4+o5EPN2hMh8iTrpqJ9Kl69ijn4bMQKRwXHPBof2YLlV/b1zl78qNzmwBUMUJ3EQBL
tZ9eg92ecG3WyOKC5h/EuQYhMfn25VZcJBN21DZkgEDVOKXF/uXdj4Qnto94V5qHa3P39O1ePeEo
wICmAzRuzlCIXALAO9lGIoat5g3LMPJPsjxTgvJLFv1AeEU4F6r6btsiniBzq+QIAUyuVf7Z1kYH
gJQ4D5bOlL+mRPT24eGsoDcfRJyV1l7SWBUWtGWBO0uxbLrCDJI3th289CBXXfyztfQiypFuuQqF
XAx2V3rBVVuBObtESuDmPKCaF+sddOa53Wb5iiap/RQws6NhKDfOFFz4OsIokxcUXlIgfZwHMd54
e96dh5ttoXGdeVaCm9gSxdvps9ZMobPydbyAEhQJqsO8HviBsUQH+ZAtuoC+0GDAgZxzEvP1H3fk
qqGddsLd14GjtS7cde19pVeYStbxH03EKdmi+hxjwGNOpP9XWkEiJgiYar6gz2h3t6pEJeFAP5v5
w/dqBaqmXOJlqMaSYmH/t7nTOkYkTANYS3RTlVN7NesjWH7L3bAm20wjtK+Z24lq9ZspyJZjIKTK
Kia0VxjFsh4PoN/fiW6mZmqEszd0CD5Ymw7VvaocyYVB0Uoz4j7QxQCkWdrvl3vKtWzRnP64r0/v
weSUwCPLJVwoUH3XaZBAMqTA+Pc54aHGWDoIkT2Ye9VxRgffJF/KC3Be3xlfTlZAA22yHpxiPU58
Mw+89cY1RnJH6VjdNqZbHqYNxYXFdHOp9teEDxBqZ5jmkFV3vFEbSzAH7K4QRCi2zlEZlBNVWG+J
igiwaBZ1USuMq5KxesmXi8vUmb8XecxWghopnNIxcm2d2eA8e/gyKzXvIryjpgdJyz4J2VU9Jydn
5ecKQvY7CArKsJkI78ifUpfP2ETC/moTZiHemv4IxE6GDTRPOl4SCf3NaEDFEvV2/4Bxv+0g2HNG
ZMMXbOE6Xq8lD8wb7rd/bn0QS1NZi9tnUjteNHFbTqlkOif6mdFlJQURt5RlU+kguII1j0DVjDGr
baPzQmuEcnEaAj4mHtxsQMLH5n99xCqx92/I8v3H2HjoXcnL5BiSGp/3ZKrQHTobVBqBIBukHqdc
jJipAOU6zcwcgDRrYi5GwvcqrJ2YxJ+l+wSvUfaOedG1BbpVXRRewpozXIkbv5vBDhDPjcCfOCkv
42+TCWORMsOOs/gwdOh6TLMm8Muy/BEnVFAuFgya1M92BFW2tBdpjEoGlo71QXfo5Vi/u+NK+6jJ
Xz3pmAoCXsqpnOcLCWSuTV6XINwq3cSka1FjgSzfTS3uFwMtzomL8vvlTigKqj6N9RhW4UIfTSuW
2LwAayY6wgaxmoAwrb9O1Ai0ErrzmKbJbI4qFfBnrNE/YiPOrY3jqSw2eoDA8jAWZUUSWy5iEH3d
WMml6SZewOuFrpqmpKr2oWCiLfjBTDgbjaaYt5fwK83rNPu6RIQkX6ZGpDa0MpRveaIT0yRvkU17
14E85N054RubrPVnu82xmibxFFFW2UfAt+bepKd4qTyRt+i0/dakow3YnOxIXHKV7QZXLAtu1SN9
sL+paYy3rgCN3hMHKmaNKy35NC+wpVoZgYb/HqEuvw7UzxniTwUcT4xh9N7gHJd9qLmwPm6XQpgh
RBwiSFln2fvxkSw85cInW/wkuuOLllISyuznlq/0walBdp4jqZNnn/uK87HVzjWRAUe1RWtd+SMA
37eegl6DDfyFCssEALhhni4RRLMvigFqxK5S/MYxvJlmbLQS5USmPq9sZtfICo9Q9HWGPLCDRD5E
AGr/vHeDRYwAPE3nyP8jjbBQ0LJbxH0yUkxN1vYQDL171lvCBMCOw4/AIdaqhXZMkySSP8df5tSO
Wkqa7v+Y7rKKc0pmWSSisVBY8Zp6e8Vydd9HDA+0Vaj4T8nKP+7ch/vUakMJSKJpEMJ0SJR6ZP0l
pn/xPH1/A93k4+aMgA4//XN+MNJ+kbVFCZe53FJldRWmLC/WG2yfV+lKZfIoK+DKLI427GYbdqoH
wlfpZ2LEUm6uQjheJ5wSQ0rpoxv+6R9rgGqz4KXQOkMgZnqA1L7qFtYzvCO0JthHPzUl82pogwy+
j7tkNbClaH8DjOYyXFPmVxzCi3ASiaatkco0g+JDUyqz8RAcspvQTLJEv7Dgyhrx2OS/OHDqjYAd
aXEWeM79IaWYuowMWbL4cI+X1Zd12vSWQj6w9/ZNNixgCXQJV7uFV6b6Rb9SR9eNKvbYxVW5eVaa
xRcqp+Tl6keIp1GLNp5ewEkTA6Xwse/4revnurit+elj5J6+gaSlEoo8J6DffbHvSPqjSlSPFlao
NL6K/k3HDgZCi0XatE9Kxrmmv51Qa5jwF2Mby9GLz/L6KuJ/k3snq+JWxRTe2XsPascgQgqx6u2w
6yDnoyxLmw2Wof65nWHp50lL1y51d7yLIPg3miaZRaupIJP34kH6qKwIdaWkGX7l0AzBruoxjDKp
xNmr/P9Elg9o1pL+haDpKIjRwz+JW5t1R+DOErvq2BfkFOtbKi+VArKfl1uJSlBXigAyB4IARpsi
9XXuaUcbGbW0fW5qOfpvdKDABm/fodmgMttarmBJf+xug2LOQG6kbB1JeR4Me+ZEY1JIOAo79aab
BMATmtV6ZcQ2Lw1ClEOXgBXCBgrCcYhV4z5dCww5LKVSJyy2RTQ7OsyAA9Y/Ld78LhL9umPO3G5P
Vp1dgkVdYH6tAoWOMn8tbPRfFvuM4W6aAJvFb7TNqsrd53UUL4Nz53siiJHxaR/iuI3ch+/K9FTN
IGcI9gAZJDa8ZQjlbM9MVmDK0zvtHey0MyG6W2GoyeDzfBaSGiEFskSGztTc/mDYhJau0TVJyfwE
mV8VlUUpCcSX2BZsYkI+WThiPf9KrbdEZqe+M1Iw6nF6JI+Pz0KNwL1gl2ffBRWlWctG6mAlwem5
cWhc7o4uzdiXJrx/YEwOjRWh4pHYex4XHAGcAFO5TokwsUKLze2v/mCRbfCCQQBGllpchc3gl5Oj
n7uLvgbU7TdaP8vFiAs48HgwMHrsDsPOoSrPAbth3c0kOZllCciDj+Kwas71nA16lNfVa5qmG3T6
k6amMICRyNTHf+x5VR5wTXRSylkhpOBxUE79IfMYhhxCPM3dG4rrNN8MyMlWEYgwxBQxWDEND8u8
ZibfxZyRpLuiZHSvAomsrcKmdHOveLYr9vwYKu9aTKw8Nb9zxEDZutwRvxxxirFkE+/3AWRKMGXG
X1qFJdBzPReTSPeCbgHvG05OExHPFgL+s/WIIPIrbreK5T/exS7QAcqqNdwmJNZpS8coW7kMY+/c
HmPD19+gTRl4tSIXzFwDy2wTfBNrmEiNf/HEWwOxHEScijo+o0H26zudlJ9IhCHUY3e23T2uKF24
4eYddlEWPg/ps3xBuECQcZ5mRu7l40Ke1EUfcly1ENNnSNtZqzZQZNlEu4aG+r4d13/jj9qLo3eR
6aSQx/QGYclzkIKIixCYk7eXxqVJpVyiTqlV7TEbRLc4jaCEE+vdkEHaJob2R8a2QmmxhLE/Z5gS
TkV9sWOeICb1FWP58ynecMgt4z/dRYdgMrzWCdYGS4Ql1pMwWo+GGmUx5extr3CT75wywtLKXH9r
T+1ugJyqWYjIl4UmglJaxoVD3TBJDhWpbOOjWn9pLFQXq5ru40Lkc3QGnUUUmaExZwGRBUXu5Jet
CuCAHS4FqM2Akf9mcTPGmFniS4C34py/aze/6rUjPmrGlCwNzxbqb/P6ykHKZR6ggBGfr8WbeViC
KwlEbLGu9AWOB41BWjzfrbbrZxVnfYauhJcaBkruNBAvoPL+JVdaH8p08ruXar6zfQQDhNJ0mDUc
akWF1JSKCE446HELFg8WNyDtHL2yr3zxMQqNTRfkmYvhfnwNWjIeeP8Xy6Xhw+T9+AZdkYK6lt+c
lCWyAVVUIruqbjiOuVgJswayDjxvUKJyhcLBl34bkYRNjehwyRdw/RPHTEBQAJAlazCSAcwWMzdI
sc08nRf5suKmXlvdNukq8gWJXiPgztJxuxAIc8KfeFtkDLdBVEh4gW+1yigNPIbss9Kd1QIZUht+
i0CRaUPHx4f2WQIiqYPFyT6zCIO1MsrwAmW9eRDquXn10EMCV4WhAFL+0YXuIe1BQnIfaEX9PLDM
boMT/GtgfJVIZ3MlzWqwpdKohTJBkw2Sfr82wavbdx8JvnPBCalZJtycARnIetzPWppVrC+TiPyD
50GiVOz4aLXJUTvqogADyOTB5C8Ny3tMEk14MeLvoeZePGEu60WSzQ7rQ3e4FVUAHEeJoByv0BXd
7fCKp0aoXwBjSN8ZtXpGIunJfxO9D4Hna0IP2AMVFe+9sKMy4lG4SwR2Qg3zcMUZBG8s6g8AkObT
cMpFYUl4lasPko80iBSaL0jVu4sNKv/xXXbSik+1OFgvZz0GtKEfGsdLGVP0bG3VoaqXAElL3XSj
nuwy05n+Nsnz0cZ0JGh8yROZKdwl4sFKW7SIIWPmoDAzrndGK4SRKTwX5LFaNr2uB5jV2LHs5HFp
J7hSuYEO4UPLIHAu20/sK8sZ+SKapMfmljZfXLar4DOdxB9fJMW+cm6UOFIaZC32yLvA8ZmGWpxa
J4ScXAkpDjH8d0hyp4pp8HTy4rlN1sY45UPfkC3ebLXkFrcgVkvjdALpKVvz/ox+waa8eQ93RT2B
og5zaxmmWQzKQNBTN9wFJpUwMOFbdGa3VAgw/t6k6skVu7vCkgo9eNC8EdD1vuh3gVP+EH9BN74R
IN0O/WArRtwuLVLAp2YQoePMK6LwgliZMykZ7kO6oRG0uxLU6PeFWPYjonod+LZGCRhypl8UH6/H
fKpmlRDN9lfLIOcGiZ87pTpBjRbPzn8v8y3Fvd3371v1szW/kBlGHbTeVS1TRoa4/OVTsUlYyHnY
1g6e3tkUpBzGtj1KOU72zrgP/+Gt/SNKYyPnmLUdWCeN9QpHZRRp+V0r6+I3q9KMKhBbIqAoyyA/
tSnH10nf+agtEg33f+1E9xzzVYbtpTi4JT43twQfqqlDes+cOZ+NjEZWQwzLla3swCbauU4ZD6hl
JirWu8HNJySxyGYBcFixMANLeIPJMFkCcvR0V7cqlbvk5mDOyCT2E8KdW/vLF69oytq9J1sSvgQ1
1/hYmA6YtgjD3H3r5zP67G6JD6E9P4UHfxQq4BbDLCYkGRYy6Qav6uZTSblYkl5YMDAFNuBzi559
GuBwZJ7Hvz8FSNHV5J5kWiBkQ3a4EL7kZNSjv9LswZ59gbLEArW8CwCTI56Y7gHjwo02AztS/k9Z
mmXDX//nTcFQOoogg8pOjxm7ZI2BuewAJRSXe5o0/7wHWBrLhf5N/8nDNDVp0rUVIlQjR1Mb+Q8L
qrzV6FZ1zFDHeYIiyQ261jg4kC+Bsatj3w9S7OIFBqsOFi6KSZ9V3L1lJ253TCaBEt0IgUkjTT9A
kwaJ8en/hN2BBMRdrqmokgFpkojlQloWEnbs2qJLoMVqzcTLjMozDf39G8kfspiYAL97lEtprl3u
+CVMQy6be4RBTOwL+VnSqULKe3fOHQS+ZO9qFXzvtn2fpdiSgY8jh9Wjd39DdWCT0AGn3wntN6IF
mmeo/gIwlMWvczHA4cVgqGC+1OeO8WiB6ISfvNA/rdx395l5DpP5jxqhmkM3Ciqe7OSYyS7Zv9mN
zGmjdeM8BxoPTRvsTYvGn9OLwfoZAylBGfrwuwroKZOqCDdrkCo72DIm426Q90NEFVTWpLvoittd
0B4hcB4k/qyTcN95TTsjgwFx3jNXael7No073Nv5CTw7FO5M00B7FyCubusHPqqYst0+5Bi7OO1Z
ujQ3MERJvbeNOqDFKy33eCZHZVLpyKdVIOPgNtM03E22eq97BFNU3wsz4nLVK1/MxlM4FLx0fpwi
DnVyQWYqQ8nrT+TyRVIW35IxHBWa0N5EQ59zAXcdC63BEclpT1aOgh5F22F3W02oXFiFxO4rGs3x
0BzLbsnMflrDqOZEMhPFbxmPX/+Dxv/unoUTy9cUk+cXFfB8mi/130MAcrwgMjNXj71kkpFJo8jN
wGVQs2j6kvKCm0wAtPZ1kHsrNohIl/s/YZwbdtuax6y8IpJXhhgJvRj14V+xRr/hGNzjOe/7c+l9
kBk9lfGFZcTxwWV0kivrd4j18EQBZrE9mpb13YG/jLOgb03i5x5z875A9pV8wqz89qAgeXe7waC8
jY6PhASs6SO0rbPujM/t3gpYBjJ+Zobjcd+vJOqg5UDM8jOQJbmrPGQ5FAZKwB31wvBl6tAOrGeb
rSvT+vEvAYy5RZg40n2zPNwXYXXpeVICmYHRSow+Pm7NOBLGhsJsQnXm3hHyc6L7oXs95PA7Udwu
pvtifooBXQgONIUdVp2lqGUrYIVEtUa11i8BjktCxqP/SOOUmg1CHZOw6p+vzOBQt0WeJwIZMRvR
JCo+aHyZSNnZwqmLTstEGECecGgOkzqNh6ltFxY0ZWyuUW1IK88tP+fUYKvEuTJ7W3eug0O5SzlP
rq+lVVi7StJnLDJN9pmTWhSdyd+l/O5I4n2ns0wqBpCxxJRPtNHsWr0+3nq+XC57dqgL6n2KVz97
u1etkAn7E7eQ9pzXE467LPj0Gsjs9qBJ3ODo14zHgjZL8PlEyJhlMHi9EV3LgT/ojGn+SW4RUi2j
FFQ8/q6TsMHGpVhnvcIJ90enTxaG++DOh/4w4qyYZ0LomDE74EvMN73ZUhsTUpUS+Yq3Hju6kjfC
sjDxPZTtkMbqdvy6bB/ijDAoet5XDULZgpVW4zompBIeBUIWuS8+MxOj+RcgboYrjXeEvTWK2igL
9zz7I3TPWPIGrZUV2AYPQg17xtvqyi8VTZ/l0etBWZrQm7SNifweYW0rgTsVd2zyalMJfZWUOwfM
4nIiXgjoMexy0wR76417mNQUBL9gOkS6iDWzAnd/UUSwlbM0kzAJTVHw7kw9dQYq/aD778uUlUjr
UyT5u3ouZDvPIa1CwM/jkR+G8E8pnUTGg0nnzS0XLJ6ahNBr3+/XPMdAzBYWMGRemeF7ktgBFun1
OiMDz07vP5zC/otwYdHnCW8qnI+NXaWxFmXaAfAqFav2Hb/aUMl9K6iLgu3cHJrLt1PL4wGpW0yl
C8rRsJlqH0vajJSBq30jlgqdKFnQkbQGywgedbW7+6yI7gXqsQvZs9DNNX1fNouBs+sFEqHLJJZH
X2df+lgO9IN66RaoeT+kuE/zWmS+FBgEiZ66cEy22Jyx8tmui17KkMUxADpSaZGDP++O2K1+749D
4i4s0T44ipipzVRU3jLeouX1E5ffOKU0ruJ8oPNF+CaBuyXG9P6LQDsGp52NUq3OvDSRQbtpuLSM
gUj2UqhRFD+esH+xXWNq3QRvgWra0oarG9lY1Zt5duBREt+rh3a4Srq0Bce+iHqvQx0izqfTq7TY
gFqdPXnPPyG9ucqiQJeuTGeILmUUTp7nrtVjNPJjV/IJmADK2vE/iL2pp5ffbLY5kO4Ur8fWas6a
IXFYLNz6hQ6Bj49Yu5KGCAJ+szLnTuU+x2WRiVMDKaQ9l4Zn4Z4H34mhjzxOYb16EFYFzPhujQsE
DEJuSUwzhi5cZy0dxK6i3FilEIEF0HbDgUm1lNcAp7Z7sOFdz+G43NfHy4OOAkYHXr4ZvciHQhCI
NolCDfJKeuOlJsGZafyuXV1Grzhr6d770gre/csxAV5oCwCNZynZ/eRy/ny9AfQVz0S5/kIAASmE
48QG7U2aSFpu/ruvNHr1VqhIWNASDzDZyLfjt+UknHArPLyA5ykOhIRR3i0US28R4TAO4SlgNn7q
Fcs21KY1SAz9iYx1MV1AwYHOQiRrJcZTGfBmwsTDGuic/z3/dT8iVoqUt7qu2SVizxepKLVxZvgT
FNAbzkmy02hOysiROj7kFs1M6h/Yu8mRZ02yEGN9OMIqTIRns2R1sBrG2bIi4Ksr0IXM5+nCEAwU
KwtoIC5adlZr0EBuTazVxq+SQgF/Pm7LmmKe4LRTbM6xED16r5zQqN44lOn5xxaKkXPVYulhSlTi
Bpt2LaexVXlqcxQ8hKDRX53djb0ZLzVgL03/4QWsHUFRVJUyT76WxN/x64en7f1+kOnGeN6Hgviu
vFfF+oB+Hfr48BkyAM/Cxqs4zMpyQ4rj8QXGYXkW9E04+3b80OpqaqaNLi1HV5g4LH1YPmdJJSvI
QYKdaMdgDf4+ArSKRJ258IVhUVUjXc5nQWgbiuAoB/7dzYyNldbZJUl3kMhZkX103e6nFqB8U9rt
Zcuyf+lQVZXkc/GW8ug0Vl5cKvCvQb+gKFrQJQcs/6wt45zCA/Vtqix29rfXwz+2ahnY6sVR93Ie
bLbV5UAsMGOI7DwJ7+JA/gEi85G6F7aOkZrR9HdiPT+uLX7i/cclOOzeJD1qlJ9EgSLmEqaOwno6
ovbFBg+YTUf/ptWwkbK9AXl1weWHDxMAnhHSWHdHsz7ER5Y9KvRBg00RVEn9Hd19CFCPp5hl3VUr
y+EfAFA0n7Rj31aZ3qFo99Zt9dLoqE0sXKPaOfPhsQYpZd6o3euuG8PWEBjbEI3Xkdqb7saTfXla
pJ6AtQMBHSILZMCoqUkU1c5ZAD9Rp3V6kSs8yPnYPWToUBCtgYRJbCnAGTh3bWm4lNfg7z5xVVge
W463VnanmcLsy1k3t5Xih5ReDWeP2Y+/o/ncw87HlTYF22IMdNaIw8UwNPFTcyzUXwBPeZo72DD6
lenpfnqbab7FxhsmCPzRkJTYsxmLQsMC0Zv9STjggtEmQ01kwbPRaN5M7ukIq1UvoM8wBb4a8GSH
1d1XQhzTvzcpEbmdswCLT160x2EP4nOak7sHmoi8vCGgChPLLv9s1h8YV4HlLiFAh8h5icEq5dAZ
3P49ymEKxJanQgSnsxHXHY3AmwyfftvTW/RHbVaFXGCLP83SKU63XQBePEZxU+sSW1D+fN4QuyuF
PCXp94FgIbGtkNoD6qxrUsznCVGzPZhdkXDF7ybu+83KCZm/GJklNCkWfV4KiwU3sY3daDuePyTD
WE2AwBW9HBcPxth1fmXVF590NLe4INDku4K0yYiEPIa0bv0FzDXmQkiM5DNWh3jUB5AFqHcWNYPw
yRVioLgkf4iTnjNbWqqX/E92A0FCQpTXS2Lio65S20ajKKsW75rrTvZFu07BT500dF5n4whooUIc
M4s2CjnzvJjXjnPMCvtbyESPak7W2LFOskesYtHQ3NoaQcyRT+mgg4rZ/QFa4zObutusQc6S3TkO
M9XKrLzoqHeXr+ZpjJvw2F9vrHfqQT39yBmRQlGxckBT6+hQ8PZEP30IooazxF2gBFJa9Igtw1+A
GWmpfzW1hHuPFrDZ4w/VF3sm1iuyjIuk7o7x9S4rTffKnLfbeIVr1GUBFHfvUWsjgSp0uBUoqTpJ
8iKKiESpwFptToUPr/YIOVmhkU8E/A8kZzAuuVRXGKL21RUUpLcI0ivLDDzlHfXcda1mO81dFDwb
fSkB9+Do4BNqO/Zu6YS0IblGgwT22NKDtP8yj9FWJC9LG6T7cOR5Q/jItmpzw2FXsRy+AFwQeTUl
FR4q+aolfnyU4sqnRRXrW6TjgMU8dTbkMCzLsC8OzWrmNUZoa+rV09/NZEjieMmJX5lVVzUNkxTy
MEpWarmAZ/ysbNQkC+T9YBnwxwVZ2VFHeN+JOhFrR1j3yuDWP32GN3ZZBB/3Hv9Tre2SKJU/UF18
Jwyb/yrayWSyrCUs6gtWoQhe3it0hj36Wfz7+mS4/jxboLwbBVkokHB+45UgGadHKg24x2L2nLl7
9O7xcCPfDdF1rD5jQ6LVQ3jwbeefNDNB/WujiJRlhe3zQac6ey5PUHrn/ltDxJE10oTnwMJTxCuC
wMz/x31u3RMoU6MYCgq2VRuQ6ONFPdv57rQm2rwQYEyFjsJSCbHzb5+vKm01B/0xLCBJ9uoI2z58
J+291Apy+cHJOq0D6HeAACtg7NYugd+XPGlmRZZwtdrN8jza0TRSPLPiTAlzuOq9Yibb/6r9S6p8
o2fWDn4Zk1pUlZhWLOdS3oDeD+Pzq8/TAmKhgPtO6eaZy5rhiSUKFNXG0dy8/0SCuX4usbsoewgD
vrTEDj49hbuBElIfMHVvD/waBlVuB/c+hIoL2AJfPFQAWOPlX2A+3x6LyHjto1151r3HzPEOPHJO
OOydfyOs1OPPSDzYV9EoAO9UZqYCWyhue0Za0fQcCEryaLRr4lhVRxI94srKQAor5wXh3R2DYUGs
Fosb7tzKMMpnjdhiG2xdyvnzXRm4otAXaJFGky8+LIPtKPSoHa5kW9MHoX5l/6vIMNY9yDZTSP5e
QTyZEfjJbec3TV8/iIo89+XoEYfnAl2C/3HkF73+tJ8f9zKUSUXs1hrIPXLjQvK46O/4wSGQyPMi
vT1zMdkT6T092e2uL8fvRThTOsE9vfiixBz6dKZecT14MWpTJ+SVmxyYxHhyMJfJmcGLuAoWm6Vl
GSJxqXMkmSfnU+Pj8c9IZnDHY/LpFsPTLt8v8yJQ6VkLaMwv6/OuqvCVSXftS3BL7zNDsU744agD
rl0kmkrH612rjc4jHAW5GSAopBMOJdmY/h+atU2TN3DPocaIDNV8+OuSNePmUXPRXPHZlUCvJ5eL
MTzCf1WPzepfGq4F8fskspHyijC0/VeuEnMEfghSFx/E91whUDlXdd7WyOlC7rZUMP3kerloaFLR
ljOkeOJD5gGU/bW6Czv0ZzRX3UqdZmHAOgh0MYoZeSnMfdXW3Ju+ofOS+HLZ5NVYO9R+cHiTCKh7
nxLMzfvWDQmNACeYr3g0IIhtZSI2pRIQgB6D8UBKzTxS/SdNOGVwXn3R+6Cd+8Vxx3KjLrCis4QZ
xGehPJv5OmCMZbs6+HhTMNDwqtoerflVjjvWesH+fvtG3fZU7yI6piB8O1dTWXXook9k+oo9B7rP
AgX8bv0LWn7l2xlpGP0WvXjE3u26Zplhw/S1992dUB7weDKYO0gSC+C9S5NSZAPop1FW1J3T4Avg
DFsnHBWyBh6SOt4HURq29JJeRm8yqIgieiOM+D6fk3miG0qBnTg8E87KePXM4d0TRPDBlRG4Da1x
we3Z4qOldFSPMsz/JYyiFGFFZayw6t5s1U09b+mDpM4vG8hC4JdoPxQ6IsN9wLw4njnYnVAHzGp0
cZ1c+Bzxk0szVrmozJuZ4MQ+93Alabaq3uB98LtFJPnUT0O7Rr62XrXVQ0InLlyMbor5pN6o4jCE
834aiQ/3Y65fSGhNTXaQ/l8rMEt0pvaE2omrFe0Iqk+DBwMrB/CxQ++WC3MXJWtRYw0kCymxJyJZ
KkZjtAsKkeM66AaFXnVFHNAXZA8YwEf5Sd3qJkC9QYAwes6O2zMaSxuqfFcxZvwNxzHCBQdKWAwj
Qr1mKlpMGJ+nzgy0JWtfpXRXEJua1GidCZssfXWEb4sVf332okmGdPioHcDTel6gb/Ym2tlAC3b/
Fb2qx0rLso++5ONERXcCnwJ9jkZA1tia4g2cavuPIg3xy+LzbcmNsRGPktFqepChffpRjfUwkx+M
s2JzrMVuOQdmBMY4iJO++yQiSQLto/pKlIw4B/cm4W0zbHyCByNvceHAH5UNN6AOxp335uY22yNW
4XuosX1tEjymNqaaKbQPwjImc/z6e0M6bAJ/PyXKi9/yestfzwdMVlnczQKLiuV/6xu6OVg7iX1X
1PIZwa9TbOrMLfb+yp/RTup5Yapt41DfJuLJWaTXoicLhnY78o2U3fRk9X7Mp6FKPnYJQUr0F8eU
7YiRqHmWuIywG/RuWSoOGa4jSQwE+yuczOLLqb6P1RR3JVzaDRKKF3IX0oFVDgvVQiD4lRzNPhBZ
wVEc/5fy1mK+5HzcmyJRAng7x8m61sDxhLf40dTeQgKbqr+OGDVBDBfphWViymjvAmQDZHWg4huQ
+4kBCLrOKrTzXRtVoWm5Kl92VqwP71YuFvgRiiNYNnn0bsFFwTJjO4N2jPi6LapVsxmle5Fbo13s
1jp+Dv8pVK7Afks+tvlH7xyq4CuLB/kyMEEwlHbs0neoKcCDZTzJZWZxH/BzcEp8z+9p0GZ3blk0
wD4j8Hxd0APYlWF4MkcfQqLTCxDy+rloYlp3AQIfuo0yHRY7ZVpPrguEyH1TtJBU1hA0Cut0Kpq9
cEvKwmjdze2sytGaFCV82dDjrKNDF3GjEMqw3hH98RC651gNcr62DPUAy9GD3W94yUrlYuDBxmXm
lM9aNpzOtH5KuGkA9gVZTYgxTVFM16NkpjLYbRgU0V4i4dO2ggYZ5a58bapvYtz1CRqG2hR50f+j
YeAEtWtIDEhOLmTBd+3yOXtekmEVz7MXMCvkBCcW0H8bm5xf3NkFM2Z9e4i37Z1PlMOfJd9ZqrYX
nTQaw9SfaxIm2l/6DmWeSOMPkrc05j9U7CCFQkllJsIh9pCIQOXXBui6c3njgAuvfiM6YBLqqCQp
7QbzgSaBFXyAcKjLU304qQkpxTBppAeVMp8tErU57I+uG3v8nW5iD2/PuOiaoC4dNJgaiCTVPVSD
DXG8tCva3HuMCZ9PtGdzgLUWvz0MCpOzlPXdI1SrcmuCjky6DCEPvI9Os4i5aVeG1rc4DZnDKDsp
tlxEplS3jHbCGjIkH34S1vgqFPrOP6tvxjPrJEgp6f4UqzJe76mQGuHnORwXN4Em1i+hpWI2Ybkx
xMSqrAhS1lFtfMeTIbTz4NZ26d67X7IIMOLiIPwoA9PILubBcm1Zkx3v55GHnhg3RKAq7sEuR6eL
+JYUaklCigz1MXfLYkHprwIlHO+kvCQ3TnmgWk2DW2J3INnMV08mfRcRphP/GtHuzxc32JxEGgcO
CzAidCPJSVeh3UOYJQJd7hCahfacFrplm4nsqI+t9he5MVlge4UAevfwEhQT6CCJOxOIctAU/Dpy
dp/6RQ/43zU8Jj5VKhRdO+8G+bjTQF+CdzhS86ztktQOJ5uwiwJ+12u/JBwHsV2CH3NxzYhVdlhg
EfxaP2vGOgzOWQLsgoLswb1VRBJVSjcGIQqgHSHV9DPSPsSWZPXerQ7ReOL+kHTtzmnitIPPyfVc
Ldf4B9CFYM2OhuqvfG2Kq2VcmDv37e0Aa4IZvs5V/OdqCQlqhz+YjM8wsUBeTPPkx8yiP+UVdfDP
DuWD3QhmcA+NY+1tNzUB9AdsRZr7ZIqaAGYS8yFNydU/RH7RRSksiS+3LN6ybNqQHXeyGSr526KO
ADGF5jaEZ6lgLSkWgE/h3cTR0axWIqFDXthnamaJQpNL9M2WBU9+zUPCNPDm8Dgcg3v5x/t3bDar
bmPU6NMN+t8RucJfVYqaUqNckPDTxQFJRDyThwle/235IdC/L6fYbmd0VBthaszh83KiMXd55bw6
61dIES2VRoizvHroG7A5eazjl+i16smrR9IyHBsVejKMOqmmWJULW+uKCOovezmLdDR7oNPGH3kh
pnCLwQ32bfu4g21LGu+LUlxXK+mwsm7c4/Yw191ULiHjJ2GeGC/0efI/P0QzbrVAvzOH/mfrMNXl
SFXnc0MGBy0hQ2INzZ/Dtn5KXS9ZC1spVQvl0N7wOzBs/HL2ClFn939O+xUSYtUsigsv2C0XpBLD
wHampsHSAHv/rMAKZ6Gckj+C6830FFNBFvqK5hYENUqqulIP6aeYaswR0F1gn33dBqecxUNM/Y0U
97UwpMuRQf+0tY0G5yz2dvXaObMPApGgxyVecAPP649WJiIXeKVssYG7UjuofHu78n7Ihs3bC6g4
ycHmV6NMGfWkWI9JL1XoCYit7eFIwAp6Rs6CaS1+px0Z76xLiAVHcJkiyrSSfY9lZF1HEqzo+iSY
hob57nDB4n27XGGJZHg9F80ILos8fdU6n733etV9YE6msajyaHzvI/rBGms2Y3567DmIY4Qe54w2
/m9AqlqWAJqkUD5Hdsjp6QH0rnIEm2KThTL3NJZ1vC7CWGEqg28imrgEj+82tUhfxmXNyQai4IAJ
NUH8xEBVwcTZ0VVM+1jHUSGU51/YOgebPBLMSAdiyAU2q27ufP8n/aPxTOb43tWQSJAUmQ9ighkm
MJWi0pbt3G0es0GPud7af733sCcA3cZcU6oaYGdX8SnU1JWAg54BzDeNbL+Jp/irl2aYGWxhMKjA
EBx3LJpp9yHgFAfWPxB//+0oF/4d6XIH/5oOjGcosTI9fwgs8x/ywrUU3AJqVhLQZTX6ATufXJvz
dvDLcNl3QqhyGxk9Ozg9I36D+8XzNXr/nAfQF6+9b7RNG+SlXCZjEJK7FBjuND+hLU/vTEyJZkIE
QSUCPhfn7K456j3cXI/RKiXWbkLF1NubcL0DQO77P5vN87R2ynezq6MHJwFjGCwWoyCrlmFMprPA
OMbqynkRKtblO2/KMyC9lx5ifhYtzdjWNpDoP1x61nHJMJmCKwar9g+0z/jC5YRFFtk6GWDUBPm4
vjo5pXSnMCOOSKRh/G92qb3zYOcET77nBDH8/qDlbjhs7B4d3f3dVVPwEHrHeqv/Edb01p9tYOad
avQwyMfjQwc9k0KOTtPWO3S3mfocP0BhBWiRl2fClID3iqRyfPU5uVBeCZx8u1aK413o/Nu88twI
3/6XqgQJUOh0HVsXZjQ48ovYPe9BxAzOKFBIdWW/rWxOaNtN7NYkJuiMIRNb+ruMMO11tjVDxMkG
QMHUs0UxVvP946LP2545Ik4oD8QovViQ01hRJAXgXhXS0haaXWI6oKNK61caIU0FWFxZnHaVzRr1
DJANAcfLl/Ky4zA/dL1ZWHsmRYRjKJuneTlAw8IO/pse2S+3ZDfB7v246oB0a9vK2CZOevayo5s3
E9uymc+YwbfJmZMwMXzww+icu3cji+7YKxsV9uRx2752tWt9sB/6Itw9+A3Y7K6xOpSfth4ZGHUZ
E/zhMVwlojLUTZxR7rpZh/wdT6uHmPUkC5i34akWu4/eJWVIWzpOTZZgMrEQQ7a46P0vemSpstW3
QUJLsxc6xNisxuvmDikn90eUn7JI2cxGDVEpLWsPfCQuctqhaK0tIB/ZVYc3pIQPFCtiFM1Tmq8Y
tvk/sOc9mO0hTGHfSQ0SY33723Z+2j/jZzhJ/KJIa7vxOdFPcD1ORUWt3e/mZW2dNf2msh9ykZky
AF/sOyptBaZn08ROiw46mFfJsHcDSpQS8tOrTnMBLWrUMQHaZIP5uJAn0YICNan4FqkJSH5QqSQK
5d92ydu8VQLviVh9+sN/Ox67AmGnqJmfv0SzcnxubDABuji/5JFi6BoXlPEhnjdGM/DFl5u0+lPL
lAnla+fJELrIrlnD8c7MlNRLMToRYbrMNtNezxuWqqw2u7cCv3Brz9nh8cyJXugekgc3JzE2BT2E
Y2gt2eMG5NBYZM7xpDhmR8JPKZ1u6Zbs8g1ypFoAn6HC4D3vScQ1q5/3sfckDOm/SyaBvtsDC+R4
S8Jbp0g5aMMGSFLO6764pP5BCOAob+OXgE88cvLc9c0cMmBqL7KcZppJzkWwSpIw3nB20r+J9dLf
/c42FI0jQObIAzjtafzp3NXMSafRsDe51JERtKpjMG3Ol9TCdRPshZV/epntH3AQQeSVeqDYn+oV
D9gk33lzrBCSbjC86qkyL0+3u4fpVu8iq/tylCXIb6ycKkQCalJN2SLulp4kRuXDcKjOitu/uPek
yPxM5Ee1VOjPevCl/rqKUPvHke6XHH1xppbgxwpKmwxV7URQJ6HvKWUZ/p/MbubLzRilvGi/ZhR0
4AfeFvTv144/D1y2fDeapI/LUoSacGAwU1smHrft9tmise3Zm+pSKFX5+YCw06pXkI/TnyvBl4/9
JgM0k8FFHcUuDk3IeKSSfbnAZ9nQoJ7tzPg0rRKLzsuE7XbOFC9y6U3aWJiH0ONFU98z07eCjUIa
JejgStmPKme/9WFgjXuuf7pMrzayNnWWEFx0EyjSQEXagWoIojWbGWawZXdejzfNd/BrdvWMh03d
mjN6itj0KcUwTZRhAbayLeCmCo7YeknET6ZFedVTeMU5dIwpP65hIa2kBOuG1ZaArNOMG7hS1Sle
6DPec/35hLdgLvzBWuCZ68a2OFn5Pl8ci/xu8ee6p9X99+ykwis9cpv8cv3F4XYFZLefPPqqwohl
JKi9Kq3nIG51CiUQ0HnKeUak/7eDR+Ejjj9tycGUTjI1jbzaq9/tZsIokDia920UzoagzVNb9Bt8
+U9RIxGIiBXyiik3Cikl/aQrklG+HXdCqgjU6hCH9lgjfyeK+SAW1md+Jeov/r5O5PJl4Of58wtT
is8YP99RlAkdrN1XKnZQ53qtNGAEvNoRUEPri7msNlB+Mcmr2YEOWKRXaYg+3VbVc2kabeSSKefE
5D1yqtMz7zMtPk9tcP5S0UuoG67yWdFYaIWgOd15sH26YzJxOa0yxoLKQLsxhM1TfiM5g5sgP0Kz
pw8gjMihJjy2qTxXWV/hHgj18QdwFCx+fu9RNLjWYiMyQhsSEvnzoOabggsN4oLMC7m6ZEloucU1
jFqzJa3XdIXWjQsRSc4pSYihc5eCCDhKfvJJZJrfdROii1uYztxzjjFp5anvFH5SJhI+J+z9stcl
HXrMmLAGNbM0U6Fc/sKCBJDjMf0Kb1Dxpx+MQJi80GQWMLVSqu9b2HUh1tHq0WMCkAe7CFoYeM8X
TFw01zXZQYgpw1e/xd+/+yiLHAU5AxbWgY0QDG8RfiSwOvlZdTCeSgLX3PGJ5nweXWnByLEy1Mgd
v75vJPiscbQH2iqDY6sM96inh0vlAdwHQcsG75qjWC8Wr/sCIt0Azpj8u7jflmIpVMpyPQ23GIas
cpBCB/Ye4Zs28RukRSmKfCc7Tx7IWunxfqf4hLuDk8iqG21J/W6NWDNoHh0MvWOJ0kj24VeaC34n
w8Yyd/cMtUica0x4PXVCJtD9mFLOk7xGXJdM/6GSZTw1eVSHl7Y+gGFBew3CLXc8r0ZXaGjwbiRu
eAn/gxB+655zFBtx3KBjk9ov1/xQ5yeeTb3AX8o6WpcdfN4W2+lG1UeagBtN3dtf+aQnXKEvtLle
8rbUtkobTMZCMXv80qZvbeW2q6nZni1EJina4iUlc4IIGlE0x/cuMMAwQ0Ss5plQD/+hLG+ia3UT
Uu33/E7UuRR/34Ijb7r9cDio2i+4txGLaOLeEaol/QHClZAgjXn9/YsfL/KPaoqs/0Tjjb4x8Q+8
3x5G0hShdDwxXe47RAWIBsO4YlVlp1f5XD5otH9n/MSaTO+HhxyGI9n4nb32hlzthtN14RdiH9wR
RLTGYsuZ1uBFnk78hNhS0awBIiMW7Jpis5Xiqniv+6cBmj0ZOfcntxHVvSOv2s9BSQCWFbbOiyHZ
1orNLhx038+zaQYeHTfknD+E5r1/VCY9orebPgayXsSaJxT7HkYfqka+mgO3LEpUTHXS46aevb/8
fKMfbG2F3gtLdLH/Fa+abNHcJgv9aIQCCvQERvZW5nfZ2CyAaPdTQDcLY6Dk8eDFTDuBUmbbgjK9
JWQpiin/A9jiHnvgF5BDSPzey7bXXOqCVIOrR3kmU5TAdGxTVuAU6/LoRYiGQ2W8RNsZhbGAZVNk
O4EiDa7D8B/Gym9lFFSqnp1PSHmotKjjcf5zFcMRnTJM/Q2UJVnaAbwub1a0rS6awpen8/kwSsmi
Qcbos6VcewKGhyJKgPCu2vATubAURif42XMz36fLc1veixsTkwvzcaoKT+ytAJ137m7PEsGlZsGA
lvazwhSIUF4ehvM9CmPgHgPVkoOQp+ml9sWJ2tEKkIeFs9t9fscBNcfdaGs6fPXSGwM0uBAOP4Km
hHhWjp7pE49D1krceKubpyyie/ncmRK73xBXnAEi4HHf+yqGvxoZKM1XGdutYX87VrFrQAsJgdOu
dneCk+8F4eTgcmQWfNKrD8ZtDF+PepZ7cBOMPNMrOvwBIDkAaXRjFZjervMXNODt5ipkIo1EHodg
7vdtzr7Iw/iK3hnC54yUSccE7hcImrPFuwPoLO56Iv4+cMkonlPQRgeMYR8PglxzXH5WBVuH4DQi
+fYiSf9j7NmzDn+QhOK+ngSIXBDSDF2owMgX34GRS/01i0FTIoxl83afhljrHEoYWrVrJXaNr4XC
fiN+2Gacrg4it6PtTdfcNGjDh9dLIKk0+kTeZzzlLPcd7D/abiLRYONSF5yplzF8jfW+sl0Puq+7
IYzpYvMZ6oRKCgoPBJh0IIJlUHGHHI94X79LTm67kuRXRri+zR8fVr8SIvI1xlAgdYbzdHgcwkg7
Yh+j8RwOZpQtqrzp5vmVFiObM96VIy/NlwLJPbTdNXAsRGcKDhVZq6KCHms3nvuhvV4DX7LXbRT4
sS9noIZk3aUWUY/rDysumWIVjj9XP4ugrUF8j3W3Z9ciWBj999NrWO9ScRIawLDv4HF1FqKn4liZ
xRaw4zNcxlbL4Xd0en73YTmP9Mj3dKdhq+kkWnKK4XbfZR8rds12f1q2VKf9iWDOiwMEnh4R6Apl
PYomD3j9geu2QFZ9ipERbXQAQWd7unc74Kj7hLp8KwjlucAGV2KzeHXeu1dfUcDRSt4WLi9rtGkv
kQzUzMIotOiApghyTRLSDl8ck7JddoFuNoduG05/LyUVNiaIzSgDN68lEVjnWJOKgpv3owcFVf3r
SvoiBs/1Lyl/0k29TuzrMxtERzF+B7zQ1sSq162PTxYSItKPryF8Z6i80ANTrEmuAhUHu3IpmCHH
5JtZrCE91ZhKNuINSOhPtev9SYQPcSfuZiDRcGGGOo7ZcbrkFwobalcDBjqCp3CQ8NyKSHB1CWwp
KVxleqhQKAC9i/6Pt/2LlRCVAfL1sR7z+Zu2HEewpnaERf2QqCNU7EiCMZiJtD0l6SZluhJog8g1
5j41wo8DC5qPBvsIPmz69yanTbjkPoEJdf2E89HLYLkD4Edv0UP3oL5JWPxuVSN7shNmmd/hn0E8
dhxU9U1GLnl+g7H2exoDTkoDW367BiarQ5A4wBDsGt5NsMipetrrQ9nNXTO//XgyZUQbFeZ5pFFb
BB+qJZ5lFWDB8UCXpxlRrWTb7eV2ON4QHkAZMmgrzGPuK4gEtXptqZrNKk+ovqak8f9Y+SxnWXEO
tZRRuwxXINF14C3biNb9N4HGzkddkhx0en7H62NTPMsIuWu815zlvcqoqt7bpS6cuk6WPCCOAgBv
kiBlYtREkkQhM3q9sMdK7a09D3HxVkPHleFrM8dzcOq/+aTRsbrseQCsDIoakzc6kxBUhYI0yrPX
l4MIhHKa0uB0fKlJifHCVbijFrHrtN1R60OjDk888KJu7/YoAcPOrocdDZxaX11u71NttmjRZcOB
+KzSgSGuHrpXoQ1lUKfEhQJLPVvgHA78VEyGSqRICybnwQYr1xPanTKJMw3MleXkNO49cF6K1ods
GC9y/BGlRR6resfY5+0i/anrSwXPD1itlz2E2PaKwxXFzqVRFjYsHj+By52I5DshguzcE4sFEx+4
R/82s9YLBPf7/MZ5+dTIJW8hwGqfv6bZKKgHajgskJdMtmDE2DjxmRrhBG1eeKet0QqoBWju+XAq
BYETSSBWPCP9hyBKhKuwAJ4b8c5FbSSwDu0RuZ1JGvW82dyoXT2qS+F3CrU8vc8PrFLSrMmUwplg
+orilAYQaNJwaCekP33OOifj+odEdQuf3aefJ713zRPkkQejZYTRRG9eHlSKqczHLCEQK+f7mJg5
xMB9Vo83irO8Zp3nKZf46JlHO4NBZLu5cHsvfFYZtO+6HwQ3zY2MFFazGqs2o0BCO6jvBR90aMC+
+M4QiwewDQwIIAvhwrN6O+yJNuMjCaTjVloed/TJaFWSfK+1adnrLtEuVk0ZEQxsQbuU4CoHXQgG
OVWlJ2v7YlqVfRFdBIGvdF0LyRp98/o5JFoKSx41WN8cjLVOtFlI9iNkYaFgD8An7MDhvw8eXTDx
Ec9RcM23HWlLloc9XWtuf4GnrYmOSGZ2aEFD4dJHIql/yr9GBqkrsY0izZf2GDwZKYWqeBG5oGTM
iAuN+JlIFW37+VJoAATzTOx1pqpgZoK/yFX2ZpItig2H+iR5k/+RtH8qeTG6aoLRVck5S9EwLW2J
tUHGijJM6JQDOF/nPIDBXwLD0BIO73AZIBWSYgFEqnYnAaML0hPOY7L8dSpdpTNuX/7POpfI63fK
lyXteWRnlNjOFmiHNg2YstvUmQ5i9YT133KGpdb1H9eLgDv82o9P93Hljq0ajhjfHTdBOK9MOcGP
1w7S8OPt2llweb6y5bBOKIRAZEEYENuo8Y+qk/I26rY/6BikVbsPJpU2+ZyyDcfQoh46Vpk47pyg
hbue0paSx98/WH+haPzAtiOQSHBs+9NXzrZRATksLRQO56KG/6HoTf1Uyq5cwgrITmKnIROdckme
bARZDYZPYtKsKhdnTNORMO1GBZ177OlJ1S4EZ3mpQtQsDzZmOBVH1nSVMQ/wTE89J9rsDxbExcWB
4e8AwpiDSVKqe5bAb6MdXgR7v86SJMKuNjJ85mGayn3nuOgiQNm7iOMga1vUJ3wI6HvrTPpUqWBM
1zKQjtbU7YtjNYfKS6fUs71cC4/pgcZjJNAYZlRvR1HVUkCu8sME7QBYVJOkdDSZWGMZfDyaMOpH
a6fzE/ArTlD74Hg/xELY4BeNop1/2H1flsuZzPU1c+pc4E1kt/kxZddofha/qWGIdIjyHD3OoMzF
y6kvG4C4UYxdW9HuOxp9wG+r4uRbYjQ5pgKXDAtMNokB5B+Sv5Oh5po4oUJxElp5raZM4IOAR0zf
CEDUIezM4MXTnCtJq9yiE0eS+jJ7DjUDZs+8o75Xyg8zKCF66CFUm7yl/qSY0Kgb+fRWAbLfZsd3
ai3bbC550a75IvUFPMFU4LQrs3bON8FXyolBpQEVnE9izzkLkK2KS0Yom5lU0+uO9LKzV3Je5k1i
W2qh6Va/SaBgYt2I79aWV3B1WpsSNO/YfkqnX4KJ6UDIB50De6nHemPUNEpiaax7w2/ksjkk7T+H
oVmA0h1L1ZAlPHD/dRLIRuOxIczI9QRRlctrAzy9yrTzGI9IYsfPkdCjuDwiMtdh4LNHewjzAM4R
qMscbNBLpZw12ZgVrH6gFtMJTQfzUvCUYodgmngzGjA7guguBB5yb6KTLs3wfTBwFA8B709sc1A+
jwnEWWVZ7lOnvWsAG/s82wDT10GQY4mCcBEnhYWNlQwrJ/x9+FV0QBgn4o99CIu0TW0rhezIdi2s
0TVwQftg0FYD6vve3NsTzMH+r5fS6qduzlXW1iAOt9gPnt3T+px3rFTH1aUFUlyBULWJhM2ZR87G
8guG6yhYGVnKJn/FUzjHjOCXarMW3HZJNNRGEiCkbO+/NLsZ3HlqzD8C/LMKweCOBnv4D/KH+Ady
sfrmQPe2CFLiFoEJwr8tmFuz9f0uN6xPALyx+7ZVnjWF5p0KCX8lWNT4xDxeemC4nv2tuZJsVlHG
FQMZ3+s4dLgkNSVc6czmxVfmhnrh/SDvx5/fMXVrxCCZiLWbof/TmcXTzWJzeJiCOeSVfc4NDS96
i+poF8+p8ZNKzbKwPpi/yAC1N0SzF3e3cJDLm72J5xFcKWLuAiiS2lZyVSuIaKtveQ3c2QYEUxI/
QW48QciuNNMtroWKAb/dhOW1IE16YMwYYXeSl/vBkviSMQcYrZ4lC7212UhhuiqLQ9nHJsXC7/w7
b+m6iY/wNxiIOI20kBC0ubi3QtTQhEkL+I1nE0M6bLkiToQbJFO5XMbuuIJ5WJuX9sdL4R8yEGgM
nHI9vhXwfRuyqF3VRC5ZGANAOghuGw7A2y5X4riifTMbxGr5+u2nn0XXrhyrTcuqAVyMFLn3m65n
lC9zw6tS56rPGssp/HHSEleyR+NRhQZ1aI95kuPQmR4tdW7USYDBQvPzQBnRQJlXWPYLN8yLFt6h
MGlheUBKitj8+uylqtUlhu6G3HXjGwOXDfHlPdEZhc76kmk+m1Xz5lEb7lLgkNqHnLgK62MghvtY
wbWZ/y5uBlatdhr85kgxCFXcisagcnHrAz4BL3aOTITntmHlGp6RTBbHhVbefWcN3T/UDh2l5fOn
p5qb18elVxlMuY9gz+VXQtydyZgYSez8Tv5WZcAz1wANvhAb1wEhjFRdOJUMiAQupVdRZwZ1LfFc
M1/h5RiFcpphNtE/jjSSdndLT6kzitW2/c3VcC/k/93X4Rw53QvY7YCcF68nM5lPJDuu/+YsPhG8
kd3Eo8Mt21ZbPz+WE0AUq5zmcKs/Yv+qy0D6CUytH7fcPCyXrAfUkYZPlhFzx/CBxmvqfdkpZOzW
fAjCbHLcBaNZct5ewKq+WBMOZBP2xtGbYgGeb7jNXsgAKgrjGjGOtBOm9FZq5UfcIw4n/911TfD+
yYe3S7bWhR+pp0MltVl4LQSOVBj1Ol6/o2GSRl8TwgpAc0Jz1xsriWptORlqJGB6mOFNyBVdFJOe
bJ9HnlQ92reW/jzfU0knJtY/0JUZfwVNMMTRcvj/XrcQzOjg60949Q2hPO1Gmri9XuuyQpZ5fAf5
yp/pYhug7bBunCcxE2GNHhS8yU8YnvDhia6rkk4IdPpRJRlJwrcpCjHTgnFl0ykJUoE5FGp2DDkC
fQeXLd97MMYZo6Pb83bKfX1Zuf57wqrWNB0YQlPpYM65Wmaw9wUSDfFwlKKFa9+sHBz4rs6+vc4E
Zll2mjJeBXkIH1XlW7PYLbpGt+AiB3GMWm6+huL8z8MTLOazMeUzOQM0dhrC7CBlK6rBcVI1m2Yc
Ib966raUxUq18BxxzrVb9xHPW78gmTGmRfytE39KXcYwi0PELTLpcnGGru65bVA4nPJLOzT5tYGe
2jtL6FMMipevMn8olS8mOn32ACAmolAfnVtS/Rwhph9c4P5bXjn7O7o81HwYqdHhr1jT9L0ylTeF
YgkldwbzafCcTSGga9hraQj02ZX1egYzHzJuTsXS1fK2NWbQdNWPOL3dgaoa/KdQniuzvBZkFzeQ
dl99tjms+/d/AW4JE43+VLLHOzuc4h/s7VGkCt5smX3VqBy1Qyd0NpLzTF0AAiO0tq1WUSN6tv3i
kvmh8n05VAFgrJxXPdfzLqLSPIoWyZGamobBgLrYmeF8hDHZwQnDI8XQytxnXp6r2jUbt4EqwrMH
Gf4LxiJYYvexSDdYC9zf9PH1/9G1f2Swyks+Je0h9ohf29hcvlENJmDQ85gWOdj8mByCWL1sHAJH
XO+C0viX7IwVDhoeiqnwYabX8bOJ9AfiPMxdWkZr23RcjI2fRObCchpOOCZJ/FloXkMSFuEziy9T
UuTooU6+HtrKNIpsyJotPWRHFsAzXOue8oETJ85Z+cOUVlLp8POLEo51Dh87yXpLRUYJweQBC66f
yiYveJIS3ltS5QGPH9+IHb9u70PAmCqa/jhblp/OsI/wUfS71T92JwZjUPvdIdycg0LwNq+nG+QQ
xPd5uUaVxIF4ZLVMzVedikZLKQ1G/aFAdDNPWIGGC9shqE9epr84aAhZ8BMNJTjQPR+WqYJ3FsbE
bYmlD+veQ/sjJVLdIHAH4iAphl764pqtoNGyuqle0cAImcj3B24LXsJ67eErWA4cOySSPRdq+JFE
2SvLPddKOJYBno4/GA6qGxgoqHgfXIPSxmwshGoKwKIMTy4X0z7OQTCSjF+zmRYMDZRk85Ieiua0
NdoVenmvsuwLCi29uq1g4yUUzXfi7VOBY5MPPMnFCLx1YdHpISfsRfxsr1x2Jlen4Yihr8L0miFR
w+r/+5paTw9OcQFmFJ/3tS3MqqjDFhOvM/6QJy7MUSgSGBzHaV4NYwp1X6vfuQRl8eZoIjqcEBu5
exByjoDPejBefvh/vC8euLATDopOe4AJOvzIsjL4onR1p+7FPvukd6TsUis16y+0sIvSxutPvf/S
niWhNA54LEnljGvG61vKzGDe4+YJqM5PYsxbyvNmGotSywFjx6sv6VTYdNpMEmZKdsbeJaTNgnrg
BnRpv2ZoypvgWap8YYX0b+jnwACJULzDI1KeZ1sj4M8N6FOlmdj1zcKAeP0gKDD7R1383hdc1fMl
D/FlIE31+fkLcZL73chloLNx2CiwhDIv7m3AeCH+DtJOBxNQlOVxmM6UdEx/YQ+D/gIolLnG56VR
Gi66PzVhXCb7hLHJaz0fy2ZXDMxxrNNLxo0Yx/VaF5optbj3u+i4wTEGGFkED/+3ydpKYKx3K72Z
Fh1Zk0G0gMwiIpOmKnm7HkN/6CSEvCmcgadWna0XbXvbNk3v7UF3gELnrEpb2hfKQ/9G4aZp+cCX
50dcBrEvuwc91n9zpe81R3iLeTdAKKBoaLM/KlYPIgVuGEgvgB5nmCo4JPwaSAI4uVdILgX7tLSX
9BBzDs6i//imfQrvlCz6voa5ZyZp5iDluEFbOS6+jlrkWmewj60sx3SRbDTg4SPCA8RL8HttdCQi
wWLaNIGK5O4ZxPw+IhEZbNZ/Hgfhz7Abqg+NXZbkFIhijYFG8upP1iSDoWV1QsYUvWAxJUcjua9S
ZGSbusyK4wjb4v/d+4wPpDXlhdywzmXJh97KjBBE1ER9fJnK8ygEghaWbi2wiWaNRQpGsNLYAN6G
0zZv9DmN/l8fzAUP3aBIDNHP7uxkHlzvhxPBVmttKHyjuI/lbbUd+U9ff2qui/jimFcTKf+CLFV1
w4JMeZa8SXKgdxZW5ROu1TTni/VqwtFUfWdekWvUK0VqO3m7H9y1tmAiuAG8N8VyMhTq139kEaPE
78FgqYzM1PwrWHfwpOI1y7JPk3xUHHDt7u03HugSa0daZ61/5BRBI/AndBY+gUwt2Tkml2E7XQK4
XRY2IiKyqGran6wMMjsRVRprGxIhe4aggMYxB0itxagfq2Vl8qAHBiP2jyxCMbZSxEd3SmaIoc4y
8nxnGm9XL2+s2EzwInwuIxsVp+D26cAfyXdhrYPzcn9tZKJmRbsLLs5iWEbo2tGWCjUWHa1TlnoB
Dr9xNVhv+dUqQO9pvOZg3aTnDbiNv3N3I5H2e7vwR05EGervdOzc7ofMN5dW85jAYjHKQqNo6MQY
Z816Z12xCauOZZWVoy4hI3J5P73FKljW9PJQ9pZ1q4by8wztRnkeH+jMw1gJuHvtZ083C/lKgzNL
C7THRMsi2YI5pqu2IH9KK2T9NqqKTmB6w4yPGxM5v81RkD5Prcq8NENBbEk8uJVIpP2TPkMBqLo4
AxZB0qilQ1ROlD7jp4TrMHw6J4XGWAMmyvf+KMhWvxzRjPQSYFTPEqi68bSlMiHy9ZERUHteoDZ7
2PtdBGzcq7qcKlZ0bbLMwPCAAgYYnDjmNtxq0OoJBEP0Kghm5qklciBld5WKGD4aAJZMCaF075FU
yovQyS0HmDJ1KzvAwj7H3E3/Ft66ETB9lekWTGD9H0bKpn6uDZ1rcKD8ya599orOczwDotvvM6Xk
F0ajfvnHsi5hP76VUIiGXfDp439jsPIHAA9bqC9nOXVYaJuqo+OyCOemt8Z3wBjKJXi8W5sc9zpo
tycxLLqHeYnt1gYVqXutxML2yudBRvmqZ98FRPI/Wn70tQuR2f+grvh7FnVXZf0IlrKbMx2lh9wc
/l+j+hYzjyLpcAnQXCtMcyVLpi0B26pVoCO98+xHxAos8tuR8sWHd4ch4xdRib2JIAvDLp5gm9fK
8pe60omftaQ9Tgb313I+N4zQN6moCvNULivRz6Bq5ydoalvUFyKdkOJuX2lr2ipgso6ShM8qu8id
Y7SBfIXvzML5PmliWA+7RhBJtGROv5S8tyjzIYDjKCEXOxRSX0/51t25ZyX5ZMITH31GiUibh2bn
/56lutjB9oO3V31sE1JT7KbN/sirWIeq99joqaU2lSPxmXKzoEtvDbbqV/+FyKmR2xJU9CWgBe9B
JddIAdVA6puQ7UlFfmvb+B6msj1aG4TwRRZnzlr5c9IdWnqIv/F60a3eheeTC5T2FLLrvIbtqpd3
ZqIfTjUOr7MlsVQPcUP+UfpQkIwW5W7JZUtZIiOOxGXTYqaQJxSqFtHUv5tTmGYtp8BEgptziky3
d93zr4jHwEHL+bVbzjPUYL5SWEhUhIwg6cIKb2tvNdRDzRcMp9WtWveKFcuiFjQ1LW9YTqD+5pOw
psQ9AvSkggpL2ohKP1adK1gEmavrhncY22YzCBglj93UNdxXhnOvCxYTUKa1LUBdqFCWaA1645ux
Std6y17k+apcaehrnZH0iQXlYd9OkilgHX0xSZ1i0qXUUlM49r232nZCubDkN0s4vOxhGKf2R0ek
tQgK7t6kGdc2HaBVHYGLTfkpriccSZxmPnvjCB/Ouw66LuTRNZAECgf1VVvW2hLLUjf21dWFhHXz
+xrS3Az6qjQ/AcWY8jv8tlppjjHTKT1qEaNx77N+IGZb4UNW+VnKCKlnOhWaIZNXI58AoBRGj82i
3kYSgk/nagj+/tqC73EZHiKyWeVx7YA4aOdFpT6F7sJfyEK83C5tfmD9Rh5GWW25qKZ6TRCTOgoM
Gfyv97ADSTQ9BSuZjIb0Xi2Go7Tr0scx0v+Jo8DZtGVIQ/eVPX9tywxtDgUkSoW1sVKa9hkMHp4A
L4MEajs5i7PF+UQGqrrH8phTUi6iXufKW2RPetroyfAntEA5FeXriS5oqLLHinknhLWjwtLwYm1L
HfUELGfIzgt4jtl+1dwamRpePmJe+qiHr7ctVHG4WwTqM+ZoSMKDzxSeFLUONz81y0xqL+nO7vEE
e3jPTwkKNtYBP3abRQgSLMO1yfkF/wVBFU98SbcifUwAdZXx2M0j1FPeRz8p/s0G0RrGIO6ByMC+
/EifDK8LfWWP3bB+JeXnNS+t7wfwSMLTEzuhKfh68YFAUUsHNsoW9FzBLu2zNEkHXLxE1nutQhNY
vYPxYFx+w7lcMl5gKp5OxGCD5hErQnMvad2g8jvXf12h0PfS3pFJOFh9Opd5vJNdXVsNBbxnZ57y
ko81iHFKMPKuHci9mEJi7ZJbUouzHms4YS03vOjnBK0i6K8wF+GNiQqA5zd1HgFD/gDFd32gO3lR
SQ3s0esi9dzTndqlEyTAT7uaRbNPeU6etvLuSgkHd8Z0hILQQLndDznPd2UfpFMSO9xOB97AKFHK
yQo9XOq3wdD5/beb5rngDwxVrvlExqP2AYuRE1qlQdMq5V9VCJ/q/USigSAZwifCVszhp97+Affz
/ew/LEBYGp4/SbasADBisnqof99ndwD24yGj/Omd6JVjhRSHwxXrkBiHoZOTC4PzTXnNX49pMjKx
ZJ3KUhWd0E8EIaAfRPQdtpWZYXLAucH9G5nFhqnWrsGhSbtrc4IpjREJshCS92NDStkQxRKFqXBt
cfMalMpmNafrgmEuoiLwGLLS0t6ElJy5dEOuVftw1ZIvZQUDr/Bm4rmPNqmBywqyiBDB7Zf2Fpzc
+DrBmI3zyKL+zjuvTAEKBDX4wRlbxfgmfjrsg8Am1WiHY/2vH1US6gVb/BcCtTceULRxSxFWvMUw
1V1H70NQ8NJzRYDhjS7ogJ9E7zzrFqlSIWYKO5GlcyiyhHAIFC2z5cj0h/c7wPy49o71JTqdeTQt
GN3xmaxwdY0HiUhNRes4DTjw8OjUaMNo8koBocAQCer49w3B7OfpsrE6M2mZ/Kyj1bbvgwzMKe75
s8LiaISlPeuxCosF5s2ynMAk/ETIpWRcWkbUddoyDA+MMiU1p5eY2jtpE4cwHRU84T+1D6wdfHZH
IsEyLbVvuEqV9Uos9vLg4i/KplTp5E6gtFbd824glrcO2i86WaLWrEsuLRcaUcU96wNVw7cgfw1p
RrCxZxo+a8A4RgJiroE6E+kCXMMyy13OSq3j1ztDMviHKB40CY8zJGawc7uGspSaz0A3JpX5qZAv
zDIzhEvahzExkwu5n2PqpcUAtfczj/cvaViqNsaYvTMlCKDhYwayl0uNWm5YHpN6HMdPRVm90VvP
QhdkylNUOr5Yk4KZpjngRjHW4NJDd4H+6sIWY4ANHHMJquQEf59N6C+aitMbZP05fwrr9o4bThyq
HwCZHSWvnBhedCxqHBaXNPdAohzShkTRKQDkqonqotMWgVf6dQtKt1NangBbyV+bHWkGV/FbiGiD
7BcUAHQNTv+j0jBWfQN16L91zfZ0/EkaoHHFoDwBupgJ+eKtM+kb3MEyKwdSwwDq1Voc5VO8JUcT
94VcF7BKk9wfXsTlEkqERy85AFEMQcAyTAz2/dkXAjP5+eS4Fj0PgIwIiYs5NAakLslvdMV1/qPg
iFpqq+cT6fnvcGFpXo3ZkqDU6rd/efGvMuMvHFRSRRCAS4aXjOwqD6Np04bXWsDGIbDSwA53TU4i
ETdrbKAUwqKiLcS/o6qbmvtuBf7OngoCvU8pxJid2crao3gEHb5am56YLsO7eIPSjJk6VQQriXPs
JwxjlyKMFQyo0I576frlwZKIdS2N9CbjM1SjLC1VxcWLtw4RuqZ75/AZw4ltmYb5tzHdHcpQmun+
REP6GogfAE8+nJGp6yx+y7rxWilS1di9rt3Hcz4j7vebKT1SKxe/BjfLT9bK4K+aK6Edw3Z+nhXE
x1WyerW65+scqlJVk/PSCvMtAyo03CGUp3zxfAb701XoRZDdXgy3kRoX0zq41SmzB7MgF1q1dIKH
uJsZz4/vo6qttJV0+FwXRXyeccGi91LuM9RbsKGKS2nqpJXkMk8QLKS3+KVZ6icp9yf21w0inwwY
r3v9sc8PtYFCdr6zlQ0UBJWFJk0dr6ooSv881URc8pwb7hVmCghkjvhRD5xVGHSGgV/Nu3F1QphW
s/6wTSQPxpFcWAJmYc61pSqgScL45wIXk+Sj0eAkkwL8hMxaZ1DoOMerNrTmsDKDAcYYYJjqjSnP
A6XnEhdSUC65/B2N+ZewzRkrhkeRG3AJDPr/X9aH0nr8CltGaBUH1LWeHoJmoFFP1VADNVUwhzQW
1Xc7pGfUcbe+O757ej+Uee+PAbEe+QFzoHKyva/04/kNK07ybl9uCDJED3SMcQB8IJCjzZOs3LZs
J/8tg6MrYue9cHEugrkg1uUSEveg4dCsRjDsJHckS2+Fy/LIFC98LXkc9qeb8hMvKu2oIDoAKnM0
iIMb4Ot7irQj2s0SKqXcKTf9rCA/pYTsBV8zN5wSRbN7Cc0bb2sAAkvzEJ5R6If0ipOjqwmqxv1m
7Srq2xR5hgL0asABfUryncPSSwhsgVhBLK5tr8J25nQQv8ycKESM5ZWvfiqmu3pAgm19xS/V+FsA
wT6kSw9ipQfUt7UR27QAeCOnCuCfbK8tiutM0CBwdK+/xytn8L92iZyFj++IdmY7fUsat5+lUpBb
rGf+fmP7pboyjP1rajg2GOEdrQCLBvNCui4DqUq0pxbL3wFO7tG2sabp4xSq7D4ZqDG1Zlusunlp
A4J1owrDwVySaOq2jiNdKV28k3c8L8pSYcq5kUyz0g6W2/UIgRpTlRLiVS7kEs5mZzsmFOY4AlXi
tfeKB/ES2Ogz+oHCEkH8f8H5VZjQAGZrRrJr1/GNwEmSTirwrpMt4U8OA7qESFf5C4fIDgCi6ZO6
VhDFTuZNt2ux4SYtzmEovNg8Og0IUTs8NsmhsP1/3wiC7W91Z/QroEIuKql/edAQHQuOCwrpmV5z
Ubqq06gSfCalodlaYHJxmOVkyiKo8WhfmEY7K6RuNhnYNg4siE5YjT/FYSL+PaNivig2hPBZYT1H
zQY3xZcMFR5CBNu0FjBgu31o+js0an47DXPSSvNhyQZz9qfyTuujbIQZFSeG0VarjD70e32hyvx5
99aFLiHLJ5MhUv/NQNi6LL3ke5iR/XKaaFUF57FAAEtomZAZipEp8MVoTGgx2mJQG3/Kp9OMpC7/
3OVdPLrX2vc/ViqF2/YzbgGXi+kM+ykO78CxhBWJ1FcbVpRP+iPVQBHOlg6AnwkWcvzhNvkJXN9n
san0Cs7NDIbtRuABgft3WLJIOKcZnpGcMTiEyBC71Z8mTawNzoxQK48L13ui9D4CT14lrxd6S6CN
G4Fa0CuxSVMjPw+pXC68KucXP1IIRHzir8bY3GYwS01RqJtHJJKwSJFwXG9j4CZKF3sMsOCjN61H
KRQ7zFg1qBu9SdYr1aSX0J83xfgPcrcwgojGJ1dLH2rmC9hLh2eNCTrAGQ6Ik3+5rCgKhs0BThkN
IHDnravEULFBegIgDNZAuLz5WWVk7bHZlkvMGSQ4Z39isEybXYK7f9MtOU7x0HcSxU26ZAJzFjob
wyO0SBpl9xXE2qokn/14EXtlmRJFjK3hrK4xhgYQ9agYEs5Ulc4HVxuRtsLJW+2TdnL4i7JjIska
LIwdCdG8Ayeg2JsLaToK0P63xePVBbc5RViryh2yhjvKSk0wXIEZ0YeZZenw32RDmVZcl52BiOjf
zP61Dk4BlmAQdBAe8A7tqOM0mcqD42y6S18IuySEzrtHUo/uGaEg05Oylpy2R/ScOBAP8COFAEia
+qseeM87jARGe3MsYBIlB0yqhlegFnUEdhBzEBCn+yTpIK6VLu6Pea7wWgYRt29fTbu89DQbOJu8
XDGzmd7y0Tre/CWIJT/D1hi80UtGb3RlfDDaEZiyiAdmV9pG0JEM7w6ZCMPLzTIK4GDwnKNJX//5
PuTAxn4tqt5Q0Oe2C85oTp4gLtYbgNpgAcwwOu0ZGsRk/gNlc5jJnnZPis2bAmse2EcWLKb8X6gZ
1Cn3cpPIDvQCTvVkhQZzrXVSnWvYdf80NbyAkhgXV+u+JMWM0zA1KIlZcTp3AvxNv4yzlW+dwNhp
+Uod5XajExwOn9T3yF1mpcQ71WXpPDnouxw9eypR3r67+XLNEP7fAyFWp3jDsoOykLp1oIY9xkCL
kNF0Vvkr82pvMGG9Vj37Gs6tNF00Y+XcCY6wHgQACHmQVOwFARun5EqwgOF6XXfT6LDtBQRQIaE6
FVq6TMup+gulHNIT0lNpRD/VGaRdvu21DAYKXEfw/7mG+ABQduKyPJI89JV1tO3wchm4kqCX5qHa
X5HyAorwSzu5tjy2yhQAP1DdfW5QKi3TpovZ3jNEawTQW1R29cuAbESxT/S36QH5+THdsn0s/C4E
M/DnxL6RFy6qhaopJ2YjHR9qHBFW5+eF6FCT6bdoRRng3le6CCOwg6/O8D/l9njl/w8V6C1mQ+RD
TYpOigxoHQtmI0VKQ1EDYXIlHEA0E9UEzb6t3Pl28196UUC8KciGPLhJr0YxOrhwQsoiqUmcKnhC
JV1Cgrx2zppneOwqtieLk6YprVAlBR9MgRCTMT9YK/HjxBMmnOsGIYbOLtRPIWPJz/BKCBSxST7Z
GGt2O+1JPCxM0DrpOn8i1VeSG3asdyLlM11PrQeEbilehZf0KKKYTQLYR+s1mJT7nmhvMI+OxubT
89LBUSnMBSmjMbDDZDqPcv0xXIZFLcrDSjf4LjBobsmvcIhzKross/sh3xTU1m0KbmvrNoKatTTm
Qy41RRDvHvAXS7GaR1KtPowCn1vt3gCFyUliz8nFzyC9nWfo97RITonJCBk8oJi7brimRzkmic12
xbIba92/BKHPvbbHvCLKRtFUyamMEAdDZUIUor3Elw4YMwQoAtCToJFFwZbYf3hJrKp7ounpfCwa
iyJapxXDPmWeEBVeq7R2/T+FKWrESmFHxYrGF2+/dawJ1B525zw8GZ0heMSN8+7mLCrUax5i+W7q
vR+hYib3CKK24Hi2OefQ2RX2AUAliGu799jhwj8IXf+FYpSmnjme9tJYk2z9PjxsdmTlHwCGJHWq
t+yl/ihUUUQaDV8j29w1ebZPbV3zEjjO1xSJcj30yklNfFwknBMbJn24ACqGI2Zfo4BHtTCDAhTn
fGzBlcM+BAI8U2eQuIBAlS6xgWlNkiIN1JRJFeZecxeYwr2Rz/2JaqfvHP8oTAXCI3bph66c5oiw
9dLhp2Z/SsUkqX23KqnWiLJxjtCkRcvH2YnZvUckStK4RfOkNP7qc2JFaEFwICeo0TgMBHybNJsF
ge0Ortw+Dt2jW9aFadpqvRJyILJ61JsLLKH+fpdwrEf7Mq/5dQiFUjRqDM5t6i6z0Uq0F7K7pGxM
HBtv5Xs3smYWSmPkoNefjhZHYRYoo1zK85Zip/t4BLcCLrzlCpsFLh2kZj7eSaMM5kt+sVAnp15j
JgmLOLsBzcfS2hz3rKuPMZGrRgRRRw2kEzkY3olQYH8DNklWJklG5CAFpgMByxehkqrxQY8iGoqk
CAja7sMd5kEJ4AOWpz6NfDd2/G6dFfTMsdaGQUO6e0DUzcVRY3R0D8b2r279Ysv8ERw6CnGznhAS
1qrBhZJNJSZJ3Aw03Rmba+j0rjFhGOybnGd+UmMdMVY5YsOVAEF5x0mbc83nAzKoocRKEuHFTzM0
L595Ov8aG8rQ0SsMFhKpSF/OByDIJ50lMuHBX5wbD8UYVmRD4XM7sSXziVoITlYW3dxOsvI+jKSE
Nygm5LvQjOs01nKAZy+H7cTtrwKvsygV7gqHtlmFtiXazprbcG+NnIW3c58B9CYq48NLI+k7YTd/
flx3sPmL8PcbVE27IDWDSrH8UvBysc1lavwCjhSe2rsEx3icWRDASlBikMCMSNM7bLinzQxK03vD
3PQqNPIjZ0XeuWWnrYWlQvA6x7FiQaZDrJidPlYAGo7jgEQJEt21k9lxFpbZglCBKDWslikcw6AJ
h2JffY/F+Ig67KkBpL5kxzW9maYT3OtWHXfQGuYSqXtudZO9csWp6btwrnbX0HmTsbOxSu72fRnb
INP1MoCJFuLcn6um6G/o7E2I3/MyD+4WrR6+vYcJqM/K0LDmxSAZwePhwAi/zMBK8qFpjEWeHJxD
uz8z4prd9qyd389IbTIOneZbWm8tUyanfZmWIjSG99ZFZKtvYWabYPP7a+NMefJ0w3hjaWH+Pwxx
n5igNXhJJFOwSInRtrWuf2sAu95bk0ZoBwdu3Rs2Ah5XEvjAvV6IctHvrJ0q9M8dc1OlyqgcGcI6
6bUW+pDjPUS+at0hPR83qIZC2POnowUgEkuIwfamGAFKpKD+MArJ0k4duH0xqdc2HPz+UqMZ0JyC
9SRk0SGwnr5IupncQoIfSRhIke6ZbKPs/yreXT0CRiaJL+adOVm/CBx9j34KJE5Au2dUATQ3eixH
HamW23ujHjJNMf9mRtJeYzagHrD3nCcaGYVa2fNUS5QH2VUrFflzo7bB5NyNC1boVs+LDOoBPB4p
+VjGMLtWwzAsbR99n7lB3hV0oSvsjkOEmCZunX6bCsbpOvStESFTzf0urz7qHbezG9u2oaAeaJ3h
LdOzG+AN6DlDOr+yeG4u8je3Ek9Ligs4G/5uyUQTv1f3EF0VjuJVHU/vXhmyoiv2LkUyTCZSnonE
JqgUCHrVOkQ2NVVBBPEFRmTXOk/t5jS2fc1E86qcBd50yFtY3amwTl1jaRLBd1tOXxptXA+w0IaR
XFSAuzmf0UdP63Y2nQ6E5IlJuCDRcSs09EqPVa29mbYJYVwR0j4l7E5NE4FvGZ7viSvVT56Flcfy
IoQvCtHPeiQ6byPJRVLnZFXvydBKvz4tOT48jyTCNAJkIrv0Gky2FpLZriGFQo0UMqJnk0em9l0F
fEnBeJ81fGvENouQ2P9pXWEik99VwWOW2o2oYtVGob+NG0qDCgv6gzEUshlN8Lgir+6LmC5PRzic
thaYxb/kMEDHoKlLFNrHwqOaU2kusp9ESgyDf3rRzZhFLKMzT4sHK89QDg3QOpqbMD/6GGBuN1nT
F7UU32qAqLa0nwPjXGpSmaPkv6LkBhd10lYmOIXkVnhA/B2GqIw+7R2c1TNUXYGamuuFsYPwXCwN
SihY89cShQxZnD9k6V4RercyQh1qXM7P2blC4I4t73ZBwkREI+53WxBEEXRmIqZvvxhcdNGgL5a4
LywfoQprBdZX2Jya/qOBi0mVumTcgJnZMXS/3Y3DYC/n/y4/hnQ1OlcrHmfT9Z7uRuvoUK/lZz4/
6B7s8UDnHQgfrA89Sj04fUXD3Zm1Xs8masrPcRbvt7nd+wg2fbN8VDAf/hrcPmNHIGrf1Oj5Bbfa
q3nKMeRAuPtM/HXdBAMkauK+bvHnJzfVRByEMynVcYp6aDggpnOImJb7Yk2FvwjqS198govwDZJh
dejytXmAqQAN5qEUuhWaBshqhaswCDLaHIgbE3jqdLliU+sAOo18xN9OgYt1xX0EYN162ikNj0dn
PMggfjB01p+prMuR9mT4I/uQ6MzynGFW82gUFHZxSX+hwkKe4fxUQQlpXQRP5ciRgyDpuLAhJuJA
Uz5urxQuwI5njaasRnsUUcctC1x/ZC19vyWnEBIgKXAbxbHJpimRc+chwzKvtWs3DPUyEllVCvAX
UImlCI2Ur0Ajh3EN4SqBxFvcXE7b8KKexnL2eu/oFeGjO07D6eDzKySlsJIzZnYtQB1jm0Zu1iml
Jf3ZhfEGvN3E6D1tBV/R/D0Glv4R7CTtJz4rEGJkDkivJU9v2DqMredInH1xzfoBUKQJ/eLOUdUH
NcxWfx5n6CsDlTibcZ/aRmTrUjpHpU26yZTx9ZjQZGuo82ph8L6PRxpb8eKxwWAb2qg5CLuAfRrm
aocSITzdx6YF7PsishWQ4B+a+9WhfrynA+ukPknppOaz27ppuq3WE00Vc6i7A2Ur0R/NTGpxbNeD
88dHyu20rpJz5BJxK3FU8uMX0OTEOCpfXp4YzN9bfzuIL+HVZ1n97mMGG4g0j81uJN6UZGz0cENY
COzXZ7ZcmUlxd31IOaYL6U/B/Ae4tDnHle8Fsz3axOGX886n5chEHR5nwf/D2G5KmnmOjwoUJ/qJ
Oun7ZS0dMdzgWV8NNhsLw5uGRNuK4jQQxNqfDm8pXnLGDXMizHMBHWUAr1zGO49R6pEBU1/qPyW6
LDq/O/GlNcN7UWH0wQrIX6plYfbJNdvnhPNdP6O98Sge16chYcOOUDmg1DvnVruRXvMmucLB9Os3
AC4KgnwovFHkR7A5ODEQ03g0HTIgi0/G29LnA7h7caDaQtp6TVpmSc0y+9GU4X76U/MxPgqNRdwS
bLQfkwURrrDAk9oGFkuChCbysXcT6lf5jAbbI+4sOVYfU4q1r3tjw5co1jxmrNoRPU2JQeoPPQtX
i6TgVHTUaTkR53yTOZe5ZaPo4F9jOARl2DEuFO0IaoF6vygFs/4t/8M1lZqcHqbsIlQZzpOoP5R+
bKZyB7qew85HBbz3xSzfPttlZ3ZpeoixuuTjPg3q8pxiUHUvcVCb92SgYwJ0fHa0URRxXoR4v+D9
z6OzbqfuESqzn+DfNd6CuAQOmquMHAgaf1LnvY5sdEP9Y0b8EKouIsQspr3Jw+Ig6GndZu3pgqHw
reokvqpoe3cACEhD2a8foV2fikM5sZDRrI3WIbcQgd9732TPCiqegzjYB2tSLI52D7S+xCgi3cg0
PG7+kx1dsSutvXfGv41JLNTFxeGEbQ20Wkl3GPQJPE6SD6AD8O0Nthv/yunmPeExub362DxoLeDj
X7TGJoGM68HGRBA+vd+H2nks3hprz11xCJdjXeWiu7UW3xrnm+wJJLHF4OWIOdx6jzQGAcURB0GM
EaBAN/kHZcVqyhVHInmNi/76aF6zbVdYT9a173O0zukB4CXUfnHFPMVQEdIp8k6WIdCs4UGCtgG8
TtWaWU9OUJADLNQo3cSaxWiEgSc/Ec3GM3XUcjxZwBBz7k65nxQFcri28PJq9Ij2d6z4iMDBIV5r
eDBf2IcuUPwSd1gFrKwrje9ej8piibL2jkVxqcQS+WEk+di3IK2a9Q9mvaevLCzF/Mu2E5CLM/mJ
/QDP/tGq0XVKSVf2RPNp/ZsgmF3IatAXn2/vpa8hdSEIKYOVODpnW5AkfFo3R3JwPtPyzZATOhuF
qni394yoY8tNJSXIA6Jm6P7kay25nxU9e/ARgIT+qqS0qKShiciF5vrkKAEaI4UxY7Eq1WLnbY0+
wkZ4wMrfYE36wIyrXVI3fcXkDgULEU5livcmEfXNnVr270eUwja4tKSZfJmwRRe1K/kZRcufBCeC
E/wCB6s0UTpQErwoUoxmhniBrzM8l11Jt7Lo3UspyXkH5G/L6xPAtDAvgL93jgP1eUikYVTRRYXX
HSpnp/af+sfNNgBSKlDYrQhtoqQ0oIk3zlrSqtrf1aNixEuUnwx8hxRNBo2VVT/twQPJADBDfdtQ
0yIIqJDCTVCfvx7y/IO36BVPeEcWbZ0t4R0ZgOqvu8roXaPx79TChply8VFvEzd8szv3frrhxVD8
eYl0xczxAqjuJDIZVERA2RgQ7Et4Ojlpc2nF3CB2xIFigeOCL6oIUQHD1UjtDAInnFJochmKznDz
v8VFQpz9iFL3ECbRc05B3hCUu7QVAUyiAUddB6PGhhus9XUF76iLNIlTsneNnUrIfmXb8GRu6yim
qQFKdGpciSxB3dQTM+m47WPkEzL/lE7yV+LP+snocbD+6yb8y0XHCth0xgSDXQxLY9W6bLftyZnb
rXW/YFfpHOPL4DwIQbfKbeuQCXNB/i9vDo+NIvZkOLgvYOZObrgDt3Q6MbIML+Q0dLehGiyCstSA
Y3mZs9E+jSMkdwUDTEvontJ5jEKeGFAb0NRcrhs8exy3ALdyA/rL6Dl7iHcarH1ASBVfnFjU53Ok
ORAH5IyaNb9ACM3K0SWHYEwPLLjAMTtmL308+nSVS2xTinNV77V+9cQ4vtBZ5tT8CA//BA6b2PlW
Iym1OCYMJbEAMjTUrCCrMQlKj+3gFs1WZ62yGUpzj5gwDm8tP9SMP/A7gJYHxtu15vUDP8ay4KED
FkAscg87x0fwc7Q+8E94ov8YMrG0UGN3YCqasFMKmn9GkWc2B1h+nif2bd47nIOvDyLnpxUSY/JJ
6UmQ4lygIjp2JYAh2mtjmJ1HaAmS7016ZbYb14HEGeUgCJInxybfeC2RER+dtN1d/NWq8G6wTB10
v+xVj/WTZAhX9VX9RSM1LMd4GGqY1j4Kzi371hg+g+a8+TIV5qmelp8E2EhpD22bpoEyfhF9siJP
2ol/+fjlE+A8ZP/ygV8DNKfOqdHHMa8c/RTRCODi5QuiZOFc9DsZsJswCM2B7fwKenWzSytEk6QO
Ve+fRhkbq5VKWTTgNxUibkkkiKU2h27mCIzmv0kIaJPoEFT/FS07Ev3FxhbKCTle0vKpIBdVSCji
WeBr9wIyQM+U4dEnzxwLw8QFbBI2PLbSCaRBFoyxB4XzGgk7MT5ctqHRiqePdcSFYQDZzHSca4oS
z2UMzCVC7tHSVcZmRsX6c6BtTVw3guJNB8av8LQ/WqNRqqE6Ab2/06sFJhFlBUATx5sS82P+bHZ0
9zF3zRfuTm2Quu9tZ17IcBmIlhlO63outPT+ZLsORTloF+ECgmJcrvvDvGsZyxKhmF8xB1WiwFKm
l22L701F74B92qd6IFqXN0TprcoDSnB8bf/Yv07hpnBt9ksctxyYHp+fLqorVUOL+V0HyB+PmhYr
lOTPuXt2/J1nTuhs0OG/Z+UpUII+rtX7EZdHnTHwn1RD1SpSrU5xC6daDVEaFDDf68k8eokYUjCG
rYbwFgcclExHjsKPy6BBxIi/4x4WtMa1tQpJn1vFvCbWSpAOplEe+TX1ANFv3lJ3bFrBzz+6nVyR
1pLiGa+LrdvPGsYLKLSr3/WHvfiHrRwNOODPdpZgkaAonSHWt8/R2c2VTyd31SO4Du/mgIleaZnV
VVc/gC9sGXwUA0T+KCZZK26+hSzf/j9fr+LVs8dFcz397Fb1+A17JOFRZ4hrfxOMcbyKiYTW5dmd
76qdSFcA9p0lDzmYjEedNaaKSYDJg39BHhoCYuNjW9/YHqCMhpOueLrNHkaw5JOUO+Zsod/h1L78
kVpNNuUyeIA7x6o77SJUBjxI58hgGJl6x6385/Mg7FkJ8mD4dvHdkuBGRJ5q4CUfg/OlRtIr0XLn
YL04AP//WOSvaUnbihghiRXuPbviQRT7wmG32TPZEdLLMGgRuc2W6jPqaR7FvjWr8/Xjgtuw/xG5
HkyRvGSVEJ2ziNOp1ps29VyxbcA7+uZmV/Mcq5bJiYq0pmfjyPdYvmyOzo0O8aecqKZMGlMBB48+
zr3SfOujMVrTfz4Ai6gNgtXLY/Ys4+EUl7JvHoi/LfpdYgjUXlEJNXiZtWdDmhUvHV8nEHurTITK
KL7c9GeNDbRcdRItuhBZg58rDLKJpPAi6dU9lepkeBXA5PnuKqtGqi7Pk5R+49QlZYrcAJ5tCufw
KvYdvvtob7sSM2QUD1ccZLAh+5NtCPZFhS14QyBzU4nbcwxuPACosbxeYuGB0QFpU30XN76i5DT0
C7N/1/GfnWNcDpUb9Y05JzgsqJnfUeN/cmUfVDzKuAMhjnGbkBC91fbby0nf3oXRUOIsn6PD9+wQ
MnXM1YQNyp9E8tf9375iwxcjgdq4GG//X0jp109+P5anCA2UW4qkRmnW0dqIRrFk70lWEed5UDqV
2SqLI1Bq5S0HHm0vCI63T1bUopRpuB9qjARy3Va+L1UBNVzBFffE0KkUxjxVxHl/jDzVcyGkr9q1
Qj6vsw2CRRetT6EMmmqA7BhKi+XHGtQI2FkfHDEl6EYR88qhiL6Chr+eCplUWe8WLNj1DdEuPtaU
o4NtW2CVdg8VBpLixUalTib7yqSUlVViLYNxKdjlqmVATigRUSohPEhE2HTyBnKxQIeuaJkVytEH
rI3ZRwwYcxkolBmCWak2u/UHQo40u3kqSjmSF8MRkBbu4D/hL0SshXafI1siJoVHP7JhixPirG5T
vcPEDxpuf2ADFdJ62yFyKO2FoqzNv9rbTAh8qsMBUf3iPOVJOb7t+i0VD7+EjsEjPYafMEU47Su8
28VdEwjd8cBsizzYet8EalVc/XN3/dt4cb4TJZrtTtD1dgT3laDPwXfbwNOGbd7yVtNQV5UJkI0Z
FO50vOb+RG1u/0Ya+GkWWbeiT+HuP6IDtqfqRxlFuPNi1yUVcA1+d3u2jwXEhQi0nRxHXm/O8X1o
5qM3GKseD9jpVPuHGHn3KmI2vw5ILGhZ6e+9+dKPQjZIuLxQgwr3yWRWM4xwaphrtGlYzYUw31ja
0tXovyvjhhC39BXk2AIxVZ6+UkEGAvHuVhfXnPCGY8y4/T2EJCU3hDRM7gjokJd1Rg1577EXlwau
chqF1fBPA9xUWw8dGDLQYJYa9jhe+jGLZ+IBaq4n1uQ5hBF6su2inSrjjeC+TGx4WBWrlCQMrXZw
0XtLyEsteUMu/DB153kNVWKeiJBVAXIFeh+9X+RguKJSNMr7YwKRQRlmEjtiD/QxENAquZDIteeu
kHRMlXBGk8QrTJYY9Ew7WI4GRs9ehmF5vofVI+Nl0c3sQ2fwb0ONPKKxjff5r6XCLUSv4Gj87C8f
jBJ0RKI+qMqB8VX3NbDpMOlF4vrTg4yAsGFojBUxetjhefqDzP99jcVldJdRTCIi+sZH4fMFGKea
iaVs+OLSbBhlAk+gjHO/yx+b9ZIocEy5ckZuqSfKBFnnhZXUUCL4f4vm9TdRTf/amrMkhqg0RK9x
TNDGqQtm3Nzc+uZyJDeVhsx/ecttkDZc6dk0At7WKG4/4bRnpaLSrmZiYEWENwgpNvfwNpkKGGYj
uojs6kE7Suq+j3ZVLPAnPBIA4WvDTScO8F+3OA11C0SqNGKIraFD5leBKKp9zSaY4CoqmmhmfnOJ
Av+LtLG5u8JFxsie66NV91SZFtxAsXGtdGeT3s9QDW3AeWv8DefP2kkrZZIFasJO2guUqjYN7qwO
YtQOjJ912BzCbZl6+QvXo6W1PrKaj13E9ZncY3ErP7JLCLg56VtWiJTo7arwyrZGNSlEyHdGDCtd
IaPuAzCenwmBnJw2/lFGQgfQjDRrjmPOKdSOC9i26I/dG7Ka27LnTcl92CWM4bvoZ/KBqDXD+olp
IIpdWNwSJhF2xbIm9SzCSoio/MG0+BTgyurDvUYtpIGBV2LhiO/WwqS5Q8D5Y/7ZWWoCSdWLRlNd
4ZF5OciVwM/O7OksQ5s7qAcAEAjPKFuW9tnrTWLYjj7jskbXPHhLyRAt4FlVSbYxb6Wb98dvn3NA
xFA2QXhG3VRlLId5OBlgOV8Uxwrd6j9XhzB25TbR1CPSCN4WT+6GLSbpFfJ8KPVbysy5qwWeb7xH
asVFSh/O+eG+6dA/s7g0Dm7hRxLREjfuP4jBEpJq55odLYMs3USFo2lVevOIixd3h7+XVtNljT/8
kSeADzlAjdnyI6D8SX24++Z429wQeK9qFxs/6ytiptqB3Y4P/LoEhVXqqJOV4o0ZgCE4PrP11SXG
jGX69DvDcikRByzDmgV9FThLi/+mwYftBfZv7gh+r++5A5JIlM4UWP9xuiJtFvoHYpcZnl+mtAk1
jbhaPeIhPDkF6ogkJORwIbVdtIkMU+6wwFFnoC1MukxCB9HCNSwiZ0LlPrYLuX4SKhak6wymoq1j
P2sIOt5bE2HSujg1VWFrGZnyhSXIk0OTwybYcdmWVzvNDt/n952bOYFjw1fOoUxxWI8ahv0jUePQ
Jk2h/ORnMgbw5nk6mLgim7MWr1KBsuQiNqZNVqsVXlyzBVuoK084txQap/3qNmfqhZuGjbOGyhx/
vZ326nLMaFCrZcAkyonKtM9oeWPLAjF1cwcNKyvxj1yxX1D7IMTFS9WrhEf7IWoj3Vk0070EqDUU
CnxKXs6QJYCCgDCjsOBGtoUttmjJNFwZizy1/HzxTbcJyxnjzlyU264CP9SfVLj+EB8fSwheau0t
MPJBUmdxThblCXa3IZsxaG9IJJ7gFsWGcseX5EQdZTDkUQQKPZ5bDfck9/tr+9XslMU6+cUZkv5f
dqilLNjeWWPrYeTkcuPoEzzs44bDGhF5hP1X5yk5tkFCmJfUpYtdhR8sPOwmflpsKRqxu+ghsvnW
9ve+TYnCqcFdoK6mVHdkdvuIeSzkl9TEPICGYEnNbDzaCeySntJpyUJfVBg01XvQ7EJInTxY+Xpy
XeE9Tfag+jU4cyE1LNNPHjUPmFJGGz1n57rZ9kty8ThEnVkLhyRQTSM3AH8tHiJVhHosQWoZeuX0
kZb/WGQobPFNCiLxPJ9QwoUW19VqKhfOEZLWtkUSoVdMMsy5NUuB8XVtlnC7vZaHEe8Z60MKUo3f
a0J5zTmNNkRusPpBQjgUBuvNgKQdQaZtgFKfSsNUTFQZcDwSO9Rx1lUM7jIrm+XVcKoCH+HcplUl
LR9WGxlvnOWhdo25RW7xv5JUWhFJp7/QeKOuW1g3KeGHzBWvRLm6OmDF3IlBSbw6fQMA/K53b+nT
rWG8v/gXmS/nDX6/n3Ih5HOzv2vleeN0wUzaP9MSWccCBkYkM3fhcreL7Hx8j+bP6CXwG9iSsEKq
C028VRCr/lxCrmdhAmC+nPg6f9phspwkryYX0VfodqBEr7L51tTB+a/bJau1CwwEyhk+aj5DtR5h
tDZQsppFukHliKJNFaNa9iAueL0+TYJo46TPdr/SBGCQCUxuDRty+Tg7+wAxfvFcwPkie3SsKQcM
IBgd1mSRslF3K88VR3m+UnmsvSJWAZ2lwcc3CVRA6Rp4vxZM0MOrtmZ8axpaEI/NvuH2N3EEuqVc
o+YgtLql1kupqgmGLAwdLviSNu6OpTRDi/3cfbxneidftp92VR5u+Bg9BCDbgJsWnPRMnrlv2QbP
9umPRmQzGZ0LhKCgNwVGEmX42JcFpv9EuYKlR9vfbcJ+pR5FKoHfOYVllIB7zwrBAubRGaMbZJcl
CbILXjLhWokSt5RW8ODz5PYPpCXHrapDVW07nrUfDvXMPN5D/nCs9lrLJb0o6Fub57imWC3A5KjA
jhltMRD24ZTGdTv8/KdRlc2dgUxa4GTXVNFRkJRZIMGGPevgZTjgZRLjI0TpsRFAzgRf0fZlHGas
nHcxmnYr5e/WRFZAUVeqC8nPzZLx/Jn8EhRkPJG5bCPgKnkelpsEF4YxJSkqPYlpjfHvesnhaSwK
sum3e8aibLDniJxcit6HCfYKYQ1Iee6KD5h/5ZPCk03hbIANxFdO3zXkB02Dco4U61YxDMkGN31I
Xv8GL6Q2m0Mqtd7235kleO3poIHU7AvkzBfHRzYoY3djb6s7/M9C/N5wSHfkmi4Xd5Nt3GecGIGt
ecqvTbylrBUhM1YIT+MFbBZfT3ESKZ08w14JcR8/Il2ej5gWu0scbAor7V0BTdB7VFz6b5CBoShj
En6Nn6lqA4rofKxKZWViCdJpCMubaFmc1PFKxO4s2oeNB759oetmnSQ5mtPyg0hSHLQDyd4OQ17a
5VyqiQwwv7MP0Hpj5o42gSv1wzU9KGzayCs5NX8OFcY3RSvBBLBwc83Qdlibj9GNk/9+d8s+Ul6H
jdX15Tqu7Ak7yPAOr3DO6Eph7TnoxghScvpkMJiZjTF3rAGVZ7NcM6OV68/BGdILAQQ4v9kCbsmi
gNR3iz1SXyHgEk3kbklNgb1cgSCc/oNJyIYio0D0/kx3lhoqlVc+aZnQEPsckzd5+6RlX9UqWba6
URSS135gMp4mhpUjGX6SO6NNhyIW+HCHJMCkvGm5csjuLw5sQFvOYtX1VBdjmaUQ21+oG3Zg2jyk
lqdkyoDH73EuCkf12iUf/vozXD9+OnovdjXl4YTJ6n6XDDsmTxDfPZSmhos9NlRNdtCKaGMUn5N7
GmF7D/uJSzR85+ZuQ9mesmQZVkB6tU3WJa5gCgElujNs+P+q+ZiptnuSgbRCQs/C1ogOj3YQrVRP
KV0xKoFxEK+RuTPZs1uK656YEl5y8jREJ+yYjAD9zVcsulTN/yMyVWs+iXM04XP+8QL/XwftEmVq
UdpXqq5JEuguwI+6x3ZVWeqO+dzcRbfkHa5Af8m+RocfEQi1jn5Hvh369gU7tIfgvGQZO4UDrmb6
HxM/uS1BiwMm/IgX6rDTdLYeFa0QvWbEvwsljlY8HSXj6WKpHiGc/IE0MyFIZeMI2UE/RDx/CR2h
eGIqD9djBYIuBNnuEtYs4+sWp3n7Cz18ij1YFKKNStgZNOw/MYE8QNgpkRt4vfGMuQWItvcxxwHK
bxcEojr4Opi3KuNa/0UKKX7vm3p0QQc+NdXMaGQZw1Zb7KO2PpiVoY9TVzq3nzjx51eawWTg4kWT
OHMeQJo2sxqzJB9pwDndRpB09VW9MlIJRKzqgqYWOQ468ZdFydmmg9L8dwblMFTc1xQTvaMDyrwE
yaNzM0kpAd0ItO7sj37wUzSG2ctsLqSA9yZ/ZpFyvWNeF98NClHyU1KYqltlp0eW3JbxI3KSQnmI
ntrVURWsyzm3GPzUVuGU2QYpykbvZC5HvTFoz3O6D7zHlwhhSVdhW/2iDIZTMCvUKy+QEF9AddRc
5toVoKr4bhwvUE60Zi0BWId/dfvMQslriJ/nda5VPo4bRWsaPEB5hIG4me0ULp+UWHO73k9e5pVL
04twdkL2xlZMNvGDIvvU5Hvq/h5y+y+KygsJOMejffgWv/3WA/cx/ezUPQ/6F1sjNKhzYtvnJkdD
cjyg0c6D/D/XgJdRvrvq97wPgaQTB5jUQEs1Nnm3yi9eotTyuDPhruz1hkh18PR0ulQ4H7xumJAJ
DI1WZGEDHGz1doVgky52eK96tISwwc2MiRjS4s7W4uZgKOOYDlGq1atTL6ejNDIbIUj956mO9D6x
8gXn0fwtSP5Wn4Ssig/nsv/1ubLuZ7r3cq/1n8tgXeJCt3TiNx2/Hgo4VimSJ/807lcQmGxrHpSR
YTsIL4psA/CFosrSn5Pc9qY6tgWtdLQCkHI8+WxttbxJK1eK+0p0w/lQH+iUjSva+GOX9tISIixC
kG5fmXvJCYVXgiOtxq99pv8FtvO/bjl/fOM/kIgbYCNHwrmOJZQ/fJee4LWRHLGuXj8slyUak0G2
o1cIdR2HY2++5+cdS05gqQscdyE8tvK21T+W8CUvI9fB3lsIieJJTNFqGRH4pTDZOuPN3BjbhIWU
ErD35v+ySB6n8xeX6Ksc/cdj89Cred+awQrGf9VjmEXQ9ipFyXz90KrSnUU7ub/R4xO3spYUqxZC
RzCwcP93/SeTryP5Vh0HxrFr5IwEDwEpVamUG7TufC6iX8jwHjIaxsy8jnQNuSoaoIxKfd4k8F+2
CxWSjFNKtyGMqSJIEWk4VhumOpgls2LZeEtoVa0I0XIn+vJ7y/xYpMvEO7uX1Dz6pk56NOkEKb6h
GwQY03emWt39Y83knDG/NVGVF0geDE4BiVF0HqotrHfuWILkQuRcXWJJTQZHRzghIq+L1IiLrGZf
6GYzJMh5dkYzgGJrl8lrpij95V6pYSWKa0pP+peG8aL1a+/mm2LH5wEswRtcClWX5GCMB8BamaWs
0eyp3uUSG7Tdmyz1qrUdgvZHUqrUOlWvoxlOkghLuKKIyVMsCaqG5vzuF7dm13ecP385j6JMycX2
VZGjA/HzCjnFrKDDS41gBBpAAT9vG/AqdqLrpbGyiRPlEBCYltj8uGTsg2VqiRh2lt0PZYdClkwx
lWdRyVPzaVVU5eu9EFg7JygqemUuN04DSS+oL8teEDwehsmxLg4byJE2j0XuXxZg0OECgCVXIRtx
CIcCphbZDcxJeEL2oVMm74fuLk8w6ZA9RCYHJQEv/29ocbZ2tum98AxtcIGqvBMW1Js/aRxNQoHj
rExc/LctbGA3pO1DD3HClJ68BgVmwMAYmqbC8qK4hDU4pBCPbterbEacTh5yrb+5R6fWcYldKigI
GScVFQTegjbVCWfnPVr3WE5bvli9yVdoDjLitKnQ6DDB4FLpa9N827YqMauLOPkJNSClIpbmndzg
CfyQhVDPNGYGc9+D6wrU9XZU6I1npDhA9RnKx3D2p2+EsKn0sl4mmT0Wr1rO/jQEH7MC3xAIX+kt
fstqtM+uwAJ4mweThRAQK1Yl1wBMrW3Tgbkrju6Pe/ZpNOcgqieU6uNMDiAwJEKekZPJZIa0bKov
4V62eIr/vZqdD7hPIMKlut2BESqJ7aHsOPZZ1d3I4fEeS7TsDdE3bc60YENoNS2gesRUsI4z9+wv
YnFjSBpdJJrxy5uUEZ2cCNJ2DtMyDzpCdk8QMOPZ30z/JzBzp+gjlFqnLSGCkj//1oPJL9QxFBNa
zC0YXSUuBxSti5b79+3xtdDSXWUaT6MqaLbuMrIpP/wVtZslVDfBTu9ePwBEEZvNyN6MXpFBYpSf
PqTwOXZUw2poL9eK0z/Th1BKRroQkJzhHnpTWv7sXd0FaIWkAcBOXxEOgH4ncfsrnM/ZDGOyTF5c
52BL+1+JHLhyF34Tyu27W2pGYLiiCm9Xv9LqgJYrBYJGWfwp9N/sAbWqITlVJvH/RI6lAryTrReA
114NsZPIPabbQ4Lk9oAElzV2osHW5FNaAnNaaYKIp91GmpCOyc7D5T8y2dNFE4zQgS3Wa06S/277
XajaokHIdNAPNfVwa0aiYaFJHFmU1cfzQrMn/ID6G/RWQP/aa+Z1yzHPpkF3jixITUMWgftFMmpO
EX2xDlsfeQV4diYFfbsME9VeujP7P/ia7u+6uHwYaUkNfPXx9YnK44JMX+qhHRlNZOf1JAntjjPo
UivluqwMKvZioIEXHV8YWRd2jzr5Gaqfm197TE8UABvcgu/zAJZc+v9eTlxlc0nyvjwmjE47YYI5
PEYUbZuL06rD2Lc2CABpWsgCo1z5OysCEOSANeIMkOWg58r7rG+QCIw3rg6QWilCaeVG5o0UE+n+
wjF0SU+qGQVNxXov3lPK4mMF9mRupB2YCfnjqeI4fUU7U91upvpSQ5eSk1at/isLiJBDx/ilvMHE
kE2/qv7vJS96lrdur3W87hM9T1ZTXvm7Clzy3rlWsU8ya0itubOkrlhYVfnXwcqBLtQN2E4u7Pcx
NO7mgj43NzTqUHuaklCcIKElwWAkdeyUPLdd5fI1gwGTWHjAUmyMYJ/zoIhiEQYYw5degxo1f2az
5MBAiS4SSnJBMxlJfo8lCvaWJ5+z00GbGAGdpeMuiigxz0FRzdv9uaMmXWR/T7b9ySU8h3ngUxRt
ZtZQq4pamDiJuS4MGa0emWJNuR7a6BTM9IP1+3ppKbtFL15J4N4ozj9YIEExaM+cv4JisUfrFveO
sxDjmM2MHsWaDgjfmERM7aEFaqGIYU/Bn5qLm8DdZR7DXKZ0wkFsMIbRwHVkvaFANFC6u4rx9muu
I9A0x2UtTmjArdlnxGT8exSJTPWMqeKvaT5IAFLXb8wto/fgA8HF65LTFhTiZtyIddnSa1hROh/p
frrE52g1JLmf6Ov2WJjAhcQG+LEDT5VeSKjBtkjWDTQttPMlB/9ZLyZw5iDVM34NCZsWNNojjwtU
N5ZymNDzk9BWaNAb7sFSGf6Mh8kvEso7xKlAfgkGSZXoEHdmMtns9c7jh8NtRIIFDvKPXPPDASR9
UnwDZmequ1CmGIcf129gSDOa8wxtVbUzS0AiEMRs3l3ZtCwDIbH/kdZ/7r5Yt03LxNc+HEgdj+Bg
mVvfW7nnmBR2Rwyh4FZr7thTt08lqjzzzKGWCDiYKcc8Oub3LKO2IEkmNFZrJ4tzeRIX/96D+GoJ
RBehw7rwZoGjz/GiP03LJq8wSmzt7lej9ibkkrPPIIMRiiRPAo88q/EUO+gMBX3zY7YEFwyTCVAn
OcTQJNdVKSFLxJ1DG0bbav88vztvZrc00I1DS359GTutCj6j6LEHe1fSYG2F1WoSKkuU0I3ouaLp
YBFusgTlz479Makj8fbMiBBYOJUSrVHwpn03tmHZ/xQU76Fjp+aAbA43TmExCU4s0CM4tyqlVvBg
ff+GsOrmCIHl5F/5QavE3lG0iq4SaL3Sj4cyLVlek/HYQ9hCFcDS8/Xq/1zLJNNVHURUxMFbGnd3
+CJaC47+0t8EO5bfbJMaG6xiJ7ZdYzkMJllvMydkrgetRzU1gOK93T9FMPBxUONKQMuP+nO1/s4o
kHbgOGUf+M2i1OFnvZYXNvkIJdA05sHWkjAnBWk09xwX/ZgGwCntgaNLEBrKyAKsqnS4GkInHNuG
fbMozbkRMg0tnOYLn/w8ThtV+d75QUUuBIj+c6/Bjdf502YU75aoLwVTKQh7+44wbayet7GDhJJe
JBtoFuhEdcd/1lvrUfolzDJ7Uoc5lZfql2NEXq01NqN0IPgUk5jtHPclSPT/zUr4xhJ89c1w9OkN
tpdB8v9doc1L80PITsmbGDRMjp7wzpsjPo1KdXr2n4OL/BbLLxkDpr8c1Ked7rJQAhM25xpE9HhT
QMx4nir+An4/Jwb39Xm6DtCeoo6Ie1EMwJSMa+76hmjnZaHeHLYcO3lQpDGquo0/EDa/VEp4wrl5
3g/lc4HtQuOI15De0IS2i9Sm4Asilv+kqpVDa6YLZgInsLF+SYPSH5aeW0Gn5olc4s37ImprWQLG
PI4AXtlVvB91ak0YvTie18uVeRwthZU+sWefQoFbqv2taLEyHx65PDHouRIAYc22SxlvHZba/86F
RMcYMbknlqlKzHVWxkRPNlo2z6Yl5lHeHwjQoX6r98mCG8zcI/qracTb/TJZ8KMbDemYtm+a/4u4
kTrAI7o41pTVK0JUuA9bejV4JaFnHfHH9NLmb1+BZck7/OjROZNjVEEk/AzPy6EwDLLYAWVtsFlL
8gQPenI438tfTRZWP8BvCeNMXULbbl9PPeQuirMn/rmwCGmd0DxGGSp8n6FSnPB+iKBZVKfbxKAD
LGYdNsxNX7sUhKhnGZbiWIj1lzzSWXET2iYf8Cg2n9Dcf2f4XwfnPSs9TI7u3wXE4hy1XDHLgmrf
bYZPwjGdAx3uH8IgLw5l/3E4L2aHsJTl6tgYAYaBPKGmEWRtbJOVZybCWYWjCAvDIZDrn5VGHtN1
9imQpdEgNBnPJzJS+R7ja3ovjrHVLTZ74UpQrpZUfA6ryeS2ZOP0O60IUY7DpuJqgcbK8cERL6UF
ZqQdoH84VNYffR1C2tudonlpEX3fTaWXWDXRS4Fnk5jbLOqa7MfDV4uC59O02hO2ekbWlUL+URZq
e/vOJ3Fz9BsfmNhA5MG+vGGk2AhPS/tKU0M0EbuJq3lOM34gEsjfGqaWMyOW3Q/HataaTfsCi6v6
N3i34cv+vLja3oFx3QOLF9LLcY/w4gBAuzdWqKhch3qL3ntJL0lq9APmKVdHgMSolxH07W0LKSsq
oj9NiL8/eSaW6oawaBlDoSEDU6dIep5kgUuMw2Dv1z7E/TQ88SK3XBQeDebUiRKIdmGdFCtUPjOx
xhrdttDRoKqldcHbI77tmh8hInQ6SYChFPmOl9nF2O9ghYlG3HFVTM1odMMz1di+pHHeuv4wzhjx
Tr/bkY+IWeuqeiTeZKzm6XfeEvinWbBsw75B10HfT8qnKn/DS2P5IJwziXNNQw0eEIiQYwW0dvxQ
+dA0H9V3dBLvzkSibGatqwORjFzalg1+p2og3XNqyHe9ZeXrvCr27e6Y2p53rNGJL1NkN2wE9u+R
BjQu1/SwY1S0F6j8gC1a6yaZCoYaCz7Py+LKGxr2X1FCgk3eMnAzptB4rrti4E9ayIXnG3MASpwi
FldnI74gYpHOddwSSSuFPESTmjoonyYCzm6EU4KDhC4Ff4WjvmeZ+L2AruM376L55br6Py8Ouryw
kR1Xwn1IqnPTCXyXrBUUFTl2saxKYJtScXMgNPP/uZ21e8ftAK7wgOLFMS+IUZA1ia6QGbqdmjM+
dRPoD+n2OeRnNwJC8xlnNaMqOqVkHPgnROG6PbDOzp5q/5qWROxAfBizvwCBbqRPCDph6kWdxD6d
NkX54i6oIPwlhfvbNPH4vQkJFV3j8cooauz88TEWxQVJwRyxQFWvBfyzV8eAG4gVdDd70PkE17sx
mJK6qWsN0AbHqAuFiZvzL+aYWU/LC/EwktQByrG1+yQkY4vRTT5KxBYhAzmGOKEDbr6HqZLFCHXz
PCMknd2pUincmGGHBZw4mQT/lq+oVrQLigqcvzEcpAyW6Up93agSv6JeMiA//hZpR2NMFK0s00Ex
z/ZyFIxOIviZbET6EAAMxvI8L2bYc1Xgtf7oW368aNzO4wKIwWGQmcGx0g82AK1m4iOk69iphDoJ
ipMP8Fgz+n9TSFx6PH4M5Z3H63lJdPz6t0W4ErsLEXSg2jiqmMab8GyUoMxZcMdLmUcitHZ+ZXQE
ey6G7W0f28OyUtEZaLM4BE4k7MUonM+g2tk3yEI79eeLTGJJkJEny8XhMVJCFJ6cIuVsK2mztr2c
0w+EvVomf+7vXzkcCIYLQ3crMKpC561mrCWLsqlLBaZLwJjgtlHOHbtAnbX1AU4iM3ssPbVS7HLg
d+CbTNhwWrXfpCS5+zFOmdsxYrU3KEs6PgrhedjM2LcWRBUDFyDBEJJihGCY3h5O4FmMyTf38BZv
lyM/fpwz0vt7qd6IaiHgB5hgW5MkCOcJbixK/VjO/KANDlH5cbC6gAhcnNR0vaKKzPnWuwg7YcOu
gZ0P1Qqnef+3DlxsAkdC7kqhqP9v7Unsqvlw7OSh804O+i7pC0VpsQrPdotdrw0nc0m2cl47Yfio
nKC1fqFApXpFWOnT01y557Liw/EwE4WGmIr+3/kLZk5fBU//ntoFI7ztNVqQjqZ/9a9PFLv6qunT
NEAhMIMHtSDEBk/jTGXKjUev/xwJubcJY0GwrZsj3gdp1z/V4+ohC5XtMe6/9c+xiDeA+1VjjYmG
du1NLPU6GQSTr79rJWEKvZxRdtFpX2wu2mR3APELZ+Xf4roUPH+Lgs6m1Lp3YNVAiB1f2URYQa+Q
5HT3vwJ3o8F4+DOjKOsIgveqhJeFTvRg0vw8JcrKgRF0yAw+zO8sK4OqeLCQF1RT+D5AIilUQQWR
lTgJlauS5kuwXMIPkRainS6FZRcGVu7nQ2BrP2Gtg+I4+AHiv2/xxrKZ8QYv62AIWOkDiI/ql9PN
KiLqyFOCd4he2Gkfc9Qc1rOrgz/oI29AVBIS21+fGjubOhFofpUrBVWnKVp8ACzRNE88KEc83sAF
T1deilyY4CKZZ/mZmP83sOZArv48mGYcoJTK8qxRtsa6itX4W296YfmcLPaHZoKI6VTirtu4I9+k
7wNPcIbrKdAaCvVcXsFx9BfUnqs1cx6IKIhXBSM5q9YsdPuX84m/YPTFagQqspLDta8yUOoiYZQt
9dyhKsRMfMh2Hw4MaUqB76PK9y4Zj427bPslsP7Eik7qc90o3boU8LFhXuoNVD94lOI9FzRiow8A
sV8uFBVIJPB3SNg9RLrM5Ihj5Xog9CIFcPXE3XUstxqfPKJDa5jde2mgR3EFdVmY8U69xFiBeUWD
InRsx5vzdP0kR/IJR71DJVfSIqF/dgC4VF/TZsg5xoldFw+z3PebeGbvhWvy4abdLM1gOG0tUZFX
C93FmwU6La6lPXVaNzqqRfKQ11pBL7CO+dhGH92lqnU/ta7PMmN2vPbRzhTAYVyNbA+++ZS6X0n1
apoHmZwaHU1UkLI6pxz+ztAw6wj93ey088JFEKIkalKo60YcpjkMLVNpSqbzDnkpWm2w+5dqemmu
hQtccZCsOcKLrxaKQN2Hc1YEBM+m9bvqbRG04o8L3NW6TNh7Gqcfr0UrSot2bnWG0HxuvnkKrHOM
YHMJvoF7IfQ/W1ZP8iPUiy9m04TAvck1EkWvKuNDl4h3X8HMbsG3BHux9KrGCmiA0mkeRkFsymAa
u7i6Tarh7xT/pij9wr3BtzGiCUT70jfSRROfKptuChzkkCQoDdjiSrjQT8dLtCP894arSE0SwfF3
4u6XBih1Zyo/F0BADM63KIY7jpxpYmMf9ZMd5eDs2qQPHF5U6zE80/MGnSkqHoRp/eIkFsJujJga
Gz/CCic8HF8y6mgK9xT45xwe2jWAH0Zixw/9glGMhoxkpL4xGWx66dqQAR4FOKa7CxgblHl4xlMS
KlpNzFkTyutb/5hCjd6M6JTgbczq8CBjkRTmzcQKz3tdQ2WrOHYJ+RGVQztSsx2sTWCOakO8UZMn
R8kGnOfPuq46Ro4cdhuAiF0gIs+VDwWwefMW8Ijj2klHWsdJ79WKuZNdgT2bUgpTN4O/ky4AfEUe
nQj3+E74UDBz0GrfTeVDbkF77xovCxfaeT3WHgRnUehFXyOy57hd33jto/PW1u3IAshLEqUWjAzE
OG67BVLWYPXe4/dwLGL4M45kZu2eAkbzv7g3HL2nutUMVjtJJleMxJqU5osQeQ+NClMMmKAfQJQE
Roplhjw0FFnUflbrqpoBXUBGn2cwCDPNDgWCCgIklCQHlV5JyjXpJXsu8QRkjFkDuFI24afGXtMW
cvZJngLjFznifctT2UNGDJWH2sNsONqb6Zul4k6OzrWARTW2VAgXYYx2clDOssIu521VmVB/fLA4
FposbdXH4hYlcttV0SUz80rA9aQ7IEZqOGW08QXnSixOi92jlZGzwlcG+TI+nLrmsOTmTSdVuM4G
xe42i31CoTgRniXtC1GV7MIehuFUk0ryOlokxzebgZ0u4IeylHSYVXOQ4Xvwfi5wBOQsVnjC0Epn
OTomHH1M4C2PrGWXORUINQgBzpD9koPbh9dn5D3C4bzlBP/OIHVHFAJEtD87JS2ccXrDSbxMGCqB
3uo/Ub4sp/MiL/Yj12qXY+NfsKw2co/oHkjI0S5y+NFe6bCPBUm1Y2Ntjpp2Z1S9Gr9NjgoSHpf6
H5lWxW1zz/lPQEpN7Ydd3GPCEYZ7Is3yTa8rwSRhiVL/Q7/D3dfiffvU9UKqv/t/ijSXdyKNOiQb
qPBu+eRfP5hnTM8eeOAyHYFotKQmvBziz96/mDl3Q8JfpIjqPiLEtcurSYbMv2kMgSheeUe8vgUb
jKpvVyNNNJF8jafsHjpsQpdW2As1t+38gJvoi3n5PuvwPq2SLr3sXC7en86NB3ujt/uQy4VrR+3+
YffIdW8IAqIa739/UMBfxryQlxa0OMJzVrdWRhgFBrlhk4IWcyieIrfj5YKbIOFBg7FnUtt+TSSD
6TvGdyZgACTWbRf6yOI09tYHa5metfdASHG5JRHryt8cNPxwc0OGp+ZTxvBpIS3d0ARI/o0Bq993
N46CEqppjGh9T0uPtBAcQshopqXd4FEw0ZKHc2p+NvgSzrrf+oUZ91LgT/r8iCZUaTe8U+id8kKG
MH3YdZOqeE3tAsyvDRCZHHw0b6IV+mc4lWvAVGL9ZUu3N1RFtS1vDwyZunyibp8ify2ZkSDmDISC
cXK55zTwv9zySWb7GxFW9yEMfwH1OLvdVWx2/GYKztRM0Jz/HbFTTwg8UcC+AQ0L7rGvc+6Fq+Do
aE9WLAL9G7MmHKMC57n31xEtGGUK/R8hvuYtIw7MCm+T6aq4kHUOEGjz0m7k601nPz6qOiTmT7YO
Q7xR1+v2iN0GPGFEQlmTTYGe+nuyRWUSoxmsapLOjqaR4koAcKHzNjPzgPJ7ynxET1U+3Fnjnli/
BP5o4dL3M+1q2XwgQ2rca3nzZaUSx65/xFOW9XZIlmBa8QPbvR8flPrubsp49CK3PdtmLa4e08S9
K9Upm6PotyPwHPqbR2hbWbiZMdCh1RyPLPuJazExsGmToro+Mg69ENaITIdCvgZvTb88BS1pA+Ps
CHarNFjwquEi1Ur81pYZHlrjhX39/NDND4cbqXPWKuPAtfUIsWh7UUDaQ7Gz1WMlFLIUo3hnH1Qs
X+UsWifvK7EdfngIvK+njofde9IcpezoH8C/R6xmcni4NDR1ou4amu6MlIwATqzxqUnJRFT2G8ub
tNAaU3weX0/+ROQiNIZOCarR61RXEVleqNpoWmHzSbMFKI84CTFC+09Dojkl4Z2U/zNeIK8JXdKx
LGj0b5E3ZUi8mVItFtZ8XuPss5FUjdZl/rB1cJpvbwIFX+9RUHlH/X/rcgkRPfAZ75M4sFhIvCf0
kT8tHzbiWWqyH3I7g2qW2Mr8aCqyf4g1+olcWFwy9nTiqHHur1i0dk25fH3VuIp8chWGFy94+Hr1
u/02LXft0pYg+9UXAQK4kDWM+f1O/5+V/7b+Nod5htMB6XUK8NriPmcCu/iC49j6OcqS9OMgaDB6
3P/TnR4KMnC/SyBRYlEWNDvgSoytjmzLV12lTB40ZXylolwcrOnbpzwP1SzvFdgcXfkjI2M8dF0/
mpR0X7Xxu671OtbC8hb6FkFTgSDwRRZ2Z7F/UpD6UOva/xcVvlX0e/mMhK7ZYfQukpIS4flXnCEU
N6nUf+G2jzDRJ6wAq8XWTn6ktVvH4tyxPrhzoRG7jUsP33ZmS3A2758jOI8Zk0qbfMX8uvtixyv7
/f/3zyv9eKq26+R59h+OZipRw1ELqnYLiIWNKF6kd4oHsZuJTqn7d5etH/0tfqQNApYwDLVey2bI
PQ/cILg/qoN5P1RR+foXtfxe1Qkwek0sKSdTgC0dKpNy79pK/vz3PL05Twr5nWERCJ6TTfYnjAQ9
BaicHyVhruMyAgqFUkjq//SuXPPBz+1jj8zoD1akvIkONwBixJxj0ISoosXh2bD7Km9OZOcWzeWK
80JPM7wIaqtDXx8kReOzZ83HguAr+0522RiK1dpreH1C3hAQRF5Ejd+Dy1Bz7CPHUmEyYRbRquzI
cBTWJKE46PIZ1FabtnaVo+/qaorQjOoZM0hRZzGlgI2+BqUY0PUi74LZBkgDfYu/7RpW9UlDti9S
Z5ci/3xK6e8cDEID5PLsfu/rRdLO159W5AmSD0apHCTvP4qi8y9IzhfRO2spFRCcJ0XCimu8G3Mr
l/19cli7wPIejlORZudgGRwPS/Yd2MgKpykatI5TsZXWYnMBpCzztMlHLjuPnWi2w7AB6+AJAiTL
wzPAzC0b0Jy7WfZ5ylZtykrmLojakZdkvMb2BUY75c2KGYdPA2U2JX8WtyYbnorIXwhy60xgm7v8
I2Xg+NW9MexU/n5T0YSoshV6C12/2VHBsVkHDKgYds/by1fIa85vfFz+cKgDVpoNVHJ+SI1YjuAs
Y8jjg1w4+BsF2zwgbND6nZwjCWk1pR/PxZWrwovEHGTRppbeTkhwMMkq//xe9opQx/n8YNBNTkEG
4gC8qX0zvxV93WvLFJbgCPmgVmsrmSe2ERBKqgT/wmdomTF39Bm6yJhDidMNQNW8dYq6TSQjlVW2
cBIsd8UiqT9PtLGRg9UQCOblsvCxtKTn41GhH1JAABo0pZRZzJfh4xTr86DVgB4cyjmuOBERbSHy
Ycq2ImYW/s2b8PluO7KvyQdGVT1w+u6hxpUxrJoo4B4J6R5jf7Nt6PZgFs45o2CQkfeDXEPRO5XO
FcE1jWbn8cedZtTXTWQfmjWWlQglH20XwblWHG9TF1za0Kx+6IObEDbD4840BlzRC+JndEx+HVY2
w4MUIVWoqYyPo5JGmG5TlePeUzZG++tK9QYS5xYZPoLaPXa8r6ZLVSZnAj2SoUlP/clVMngAOvyu
kv7FfB0dNDFw0vVFv8HLKktZyoZlkmnLCAve7JLR8vsn2fgUhQSe4iWof7BE1X6IU52S8hTg+M56
YwfFe+mFtNvrleAF/ciJNT3vkVbe2MW1z75mDQaOJi9U1DLiy1Tdx5KL/MeRgwGOh/wyQrOe1uUs
OegaqCsZc1RLC1HyljrdERs2b/wPpuRUzu9AA9e6l+pgMR/vcgotOgd8uQ5wWXfbEOf5vtyTqZ6/
hLIUNJqkM/IZ0e3mM5VldoqtySiY/fS9jtB/tMjuiYxpOVrU0cFijEA5piCx6ajwcVz1qVnMbUCL
P78DaQD/Q+woAMGIkFn10MVLgaddT4cxAK9rWZkh9piVgTlvQWqHr5QptzVgJtvG4fO+/hBpZ4sX
//sjJJGlQU6YMlsur0FD1dwlpqhrjVvRHRcJctsolf9dPbVA777qb8/gPU0b6tQipLHEpD+xtv/Y
o9Kzusj52L6ySvztLYVFK9PuA6FagClkQLwPfouYuGmD1oZr6x2Lm6qHAoqbXdUW1FIgrcUjUfCh
ZhYS7UVuKYK2e9Wzw9LHTKCC/OZKFINOH7ZxnrFr0RpMH0XHdRoXgFC7yrO9HjZqRTau788l+njU
8L1V2RC7b8ZXG01qBygtMiSLdfMRfTFrXzj1BbS1EInlePRwAZOLvt6HPN5+3ol5rcJzyx6VpQVJ
G+m/5yNql/pgynTwdgiWcdzoY90EDS6dNf27+QP5WFI5VvdFa1E6Bja632msXoO7hKdUcntPuUr+
meyYRJleWvr6+ZXl8Fi3b+vO2G2ASDP+3iHTYZlgBrucECxr4FR5GigsGKaHAfnmXTjIrvCK16Z5
/Yh0eCNBVIQ17gBYkuykZZyj6pjhOn9jxUH+l9d7iGdMqrK8nHc4t6O4nWVq7HQvahEROZQCF8ln
8uBh/+hU+Th2hCuvfvpCwd7uVkJGyY9IS8wrsw33gCQjbM7jlwQ+cTfQvwNQTI/K4zBUW5LpK1M+
aw0d48GtddKLJaGX1g7MuDdtOu33IKKD3NDqx9ypqZFS9i5N2iTGrgC23UHGWvesjl0eg+Qijdx1
wV9TKeApXtOd0x5So0iUncIJoJXIs5p2wxGjCGthV0UUP6yz8es51ZD8m9Z+GL9XZhXJH0tYifMv
VislUmJIIAyw7axeRif8eGFyTw3MZSJ2pvUaKLIixzqKhPvC21Nf0HXYTenTObsvDtPHH1Mt51Hf
nL92SRiRs4DkVs5PdZUdtQlq1cgeHICcG5bNGV1imaWSAiw1rqdUSsdZa0DhyThQ2OiOEYO0nYy+
Qy5Mf/bls5AfQx7GkMPeTsIQKa+1YF2xI+G3i8b+XWQn39Lk3z2bpwwhOWe8QQ4LunaxS4XN1StG
oQEFj6fOy85cMPGFm6uA3v9PUpVp4e2t4PxWmpfNnNAlNleW6JSLm0mO3R627SFDVYqybx9du0cQ
2+4d2XZaYUMHq5MckiWW7DSZ1akJORWU1i7BbKbnhYY+3l/4HNDG6CSqlfwVEoQOIQUOZovKYX37
BaWKrhgIWG+KkOY5JYTXsC3EChE+VYtjEX93UGKapNQU6+oMef6W8ux9tUTszqsjezeRK6GsRft7
5bKwdcSC+0YatB15Mz3beWTBHlyiIz4taKumPGGka9zJ/zwL1L3oTlB2MRUKrrAwBz4/J1iwQ1II
J4DhJD0dB2m8pjzCs8tp335JlQt/QFPiz5SNl20cPmPfOsEMms8ck2qvNvVwrXiK57BpfUhyTSyc
UPzDshRW+S3x9y5BMkTJbTe3/9x3+ckLKxReZQMf3dJMG+lNUk9gPlpd+FrI5dSB1IcxtAsdHuRv
baMnZtEH8VdXZ97BtmJdOWVSCCiTlfxKg82AyFX4THCpnvro+wXfRadbH3/HSpKBDljxk1OBBVCf
Z6Y1EidWhdnkfC31XeJ61gYyqyd53DU5lJ8QXWV3Ihh7wflTbtzaX2zXOvR+3eEhXM1s1qnZha8r
3p+HTz2Y6Uhv7ouPcYYvRKBAGR6AFBdC2YA2tl93fVGNP2A8kKkGGptJ5tD0OD5uIaxiZDlEMKG3
Xm4KtxaqVws2EP7MdnZ8P+EXT0UXqtuFI4fYlvtSHbiffugrE9AbuzfykUz4kJzKuAQZFZxUb8P/
RyUuh1FVOsdZD0U+ITvCODhZ5BPMs9WJRXX1qBmsqHsZorI0x8QhKqQpAvJMHZ1IpaPPttOlj+09
0MmOGQ3Gr0IhZLYU5PRRCDSlUbMVbh3MS1K2upsV/bOoZIy9l14mqnR9iEfXVI2Cn0QCrqGhpbNw
mRfcBhqwGcUcQO1fIvH8VdPduDlb63vl4maMTwmITCxCWQBitq4nuxRFCEEGLCsJizvOgsbFpMDP
z7yv8DB/1EQ4se95EcpW4IvITqhMlRYWoXoejYmC9sD3IY70uHEKkyqks3kbcKZsbAF05twf0ci1
OSqJp9K3p/Cj9DohGTLoAcbIAZ7LuZ4ryxPgOQjUaB1l0430/Jm/4hmdVqC+NjKMqKWBfRozCTrB
licamMLXUvGqBLKe0mpNXvr3hVN68Cb63YP0Et1+gewTK4cbgsvkMGEDnoy78sNhB2g3YECw2YBF
4LArSJKvzxiyWWAhKpFsvRoKKoFieVFxncNIEE16K1M0ZiTHxI4jBn9DT6H8crF8uvKhYpxZvyTd
meZQkyYgjY6E/SWRBGlmeQb0Kv7jhYV8eOUi/KUf8rFo7bVe79d9PcN2Kn1XMxdhf11iWmCLX8aj
Q5pI3qT135tD6104WsnpHf9ppJtSDubyj3nPw3KHwNkPd/OCFvEVRu8iyLulVbP4qeq3LEV0hsTP
FbhideArM+OJ65duVqguZTZxf805Yopvo36NcPVqi2+iePC2kczfWQyrp6qzu9yr9/tiVE9qHQrZ
c7vLLY1rKzX4Z3xzxkRdvcZPHXfnnrw75NYbP9ps5I4SCN36h6+TEyCjdc01zuUTrGCSFrZHgKD9
lxqr8jp6oGwPKUWbiqRCXxmhoAJqqVWWvEx5gTcAl4RqGudtCdVr6lY2qi2DqssQd70mZXoSVK/K
jdi4CVJPe5JvQyj1+/DZpl4saq6Nkmh60ong+koGBauMWB0tt8pfpCLsxzmctaaLyOS0QnQNZ4BU
k6SfkGWp8bNvUM4YLF6gEOzSwavC/ECQX+y68CJRUiPGnIshLJAkoqityrPVWms5tqpkVcD+dfw7
kno/c0W5nqYBemIs77p8Xyr4ZvApH54kITVkIvWotNL2+QPWiS7GjNpsH1tT4c4N31NOkor9u1MZ
QtOMTEeqmMa46IQtRbJZnOToQRiFVCiUPuCwO91LVaRQ3UrxapyQd9Wr20uxa5o6Xpc/hUl/k3Sa
7jIBJkd+WijLl2hB8epVHqmXnIeI/pz9xV0ZuTFddKmqYxcKzhVwYt2tlbfvr0BMLZ+CBAGOwPJg
XLxDntexO49kco2BNUwu8QraY/HCfU9HGD0p0M27U37g9T0/UxgSbOA6pvJOzF06EK7ow3f9qgBG
JBzl9y9vl1DvYeskPOrHBtsN13KuYytaSUOcc4OxWePThchd2TnxCsZZvPq3eNNKUBPAaSuBs64Q
BzHBpZJe1fhk1KCXbjQ2rAeqnk6+jBMBnAAo4xYtGouwB9nxkcpFa/j7yj1l2t+XGYtIU3wtNOaZ
/NZP2dkXLUYFwjIsxvmTmfn5x2VXjuUaDj+rNjvxfyUHuB+/XlGAOzqRv/Jjj05s/84ZRIj4GmMc
smLWxbUbVGgceBnBmznvP5aCBdmOg2yeDiLNlyvMJOcZlUWRiQ2B0NBCDyzS0cEFaOGX8eOMMQx6
FRKRFLgsTbY/oXuv1rEl3EBQx+jBF3iK+3q+5u6IHIn4LVKGa/+3jZpnXQutz1WTRKVdUogkLwnp
17irdIbqXr9k+4ia2I7XelQcZbF6aLGbSIXJ0I7j4OW8Yc5s7H/8VitM41ea212n8CriRL0sZkho
KI50xI2KqpVnRD9ge2EgwVhGbwSsyzlPjSUioNQkrJm5gMn9hfcGA42N6+E+cKL3G6TaJ4U6+91+
rr4CkfEqfRG0lcgtWyp/SMw6n+IQCNQR9pb1iYQ+Gf67G4ksGC31yJJYUaQjVVJLdXv6AKbG7xwY
wj07HvIttIBDvoQzeko01IEAUAXMOnAlKJdhJS2zIpRA+Z4BTgIs+9E+2NTR/ywgrgtCxpRX7Le/
sKZ5+404rdZQOKlZ1waNpkEjtKE6zi9iWFZE6pMf/Fpjn/uZ4VY7PbbKmyKb8zOL5SfwDRbF3M6t
IjSx4dbmnkbmU/Ly7QOjvUHoSr1HUU3znojnj08i+cztV4fhgxzQLFdfz4MJovwbygov6OTArv1D
WbnbYFKrGbUJHVIp53ZaG1cO/JQeXdvpzuy7TFgJyU4ZZ0jS159elfHqxN75L3d18VIOP+u0/vXe
LJhYsaUWXNz0ydcfc+ZZuEzNQ1fvY4xqUu+JYZnRMg5qxgdLOMHlTemHg/4fRLT4SMyllI+FYqR0
2OlPIEVu2Ho9amGGdV6+BE7lYqndhH0HRoFZwiaAfXU/l2w0xKYrpbKlTJpiBLYU2MjMNPvre2hC
+2I7acP/Ss/uUmRSo89o+8xFFK8PhZbGKUsI3cm0OAUNzoTZdZlEb/D/S1FsK5OWQm3jGOwrISVt
UpkAl+bxpmSsgRXakioeLmQV5AopZfjv34HAqkSjSv6up2kTSqObsDJwURFcjmR5qPXaMmYRpgaY
PlidIQDR9y73r2vOhJEGNu4U8x1UPrDIW2kDA5JHPUZ35Hzgbpig4m0WoCLJ37mN2+5b1RZuVfgy
jwVYRrz8W/ngScW1B1f0cFsLttmfRZ5gdn+qv4sjrHgBI6dzNZnCBZ5yDuZSDF0nWd2wOKe+i4r9
q/1Nl2UFOMYtZ19kWYZLz5s5ruz6jAjMQDB8Ikve+UmZG4s9u0m9BnDr0ZuAKDOsdVef/1+HYyfd
oTCgqUo7GxksnbEMmbt6SuvgzZeuBqaJcjgif7pAnzMxU3ME0hDMbuo4gKBnGB5g9+wmqwQsMdML
9O9+Gn0PYJuLNgxLp8qgoh79z7n3QLWkV/joE5yrQ/fA0xKnu9i7xOz1f/1R5FPVR/PwGS+UnaNc
gPqqjDxiUWR3ydPiKAFPAwc/lmuvKCVAz+zbsbfeZg+AVgt7Y4vHw8307utdnVT3yKorLBIAeQfE
ap3pqkyYTr+vicZVa+A+8MtVwO1dARndzPTBiH0xdhJHCbksbL+B+CYtUifcx9B0FTfNWu2IVnRM
zrO99Su4hU9zk0tX5sJOWbhBR2XH9B/4HhPBmtzjvpWKrndZhYNRDal0jxFYuHjhfpPUKfHH+JJO
hTvJZYW4jj/QrN7DwJ1nwK811Jtp3QIwIkDZQqhepAD81uSuga5w8dRIN+u9hlV7EYErDj2aZ4ut
0nJZ/SejI+GM8HQws0PacydYYhnEmoxu58kIJBi/llXoYFf/EIsOiBZC1E2xYWsV+IUeb+mU6jWj
s8VG66qxUFtggtrOWqLvjjnZknuHy6fl6ELz/9gwfYkBDa+98gE7fR/GjZ/jIGIHdJCp8GAxbaxI
HdtWF3dtA6Mg+wp2azBylppJ4aWSZj8GqJWO5y8MnkDwd7UKC5ydMS1HzXKtUzOHUECs/i99BPtc
MbNB0h9jrMAEuvehaxf9MTXZpaO2YczviRV1nBQAru0JCPZnOdLigF5fosvrjcDQHQvCyv68YolV
EyzyBFS4tkTGMa5U4HJZUi1Xvp1ZE8s9fzIKEtEgo/ztl5ap4inHFPDXbkAlP3C2J5Qujqoa7AcK
BDa4zQzqsyQ4WrVgXNNGg/L0f85c2+YAhcjuD6s42unltBSz3X8gsbgcu9GWFzYJnOBJW3u5gOh7
3cfCkWR+MoWP3jqBT3WC5bH98uVyBdXUXqWbAw+qu2Ov+MoHTKsUVKdii03UxieTRKRzkQr6ZFSZ
WpkvUo52HsohkUdMvF0YSAFX7m3LdGA76zqOFg0UxN5lnuIrcrMMW89oWMI0vlTm0D4vdtI7CQrX
yESddNCgfT4ndwDm+asq6S9/ajJK1trLhuouT0F/5MrzE7/rrdUQoHK5FgGWOPIUuuvYNqCXN9ux
095QutJh195eAE3lhWUm966hUnDdWQ8UdFBtZARqZCwbbGpOE7tuRcXRdNtIbypvL1+2mXdWl1uF
gDES1apP1+3f731kooycSlPLCs2kFTwr23ol5ULuvcFc73HDNnTf8ZqEW//A2v/b7XWjO6V2DdQ4
TwxiUNf0AIXI3Nf4vhLO3CFGdmtkc1ci2V8w/ruKjn2F7ArjK526U40D6UGliIS5BhPfYFNZyqtL
TyWCcrSBmd1JPB8RNUYHDZDgAqsmd9iP8Qe2hBSrqeXtKYoqwGp3kx2ndNDiTjiBhTQJsULMGbZA
FQLS4DEvuHiovEuZpN00jQ2o6M7gsJpkrIo1SM8pTxzdvmTvG6KycnqC0dZck9t5eL+MkanRlmUn
01UY04Gzpq4m14VSP5RRAeKizIBPUB4DKFB1lH36uexOcAmoLeAU8z3+BxG77IAQm2kstaTcPbZi
TFpNx36T50602DTR8pjxPGpmob1AZN8Axy5iC0sjO1SZQv+ejBSZDsD5BiPOlHW3o0qWm3R2nCax
G2Tf4f5/+m6zAmiLUbhXaXMDuZ/WoAaQYG9WgEbT3E1u9gjd7rWxoxD7rm7bjIgbidO0J0COb/e6
+d3OS3/R3gJ8VXxye1cfF0XfuVzy5kxy+QO83apt9SpYDaiCVs0Nw0N0rvWXOh0igFBI8Jqk4VU+
oXgS2lIjptPMpFjJWMjMsKdmKFUV+VV8TnKQXq575wPoo8zMQgrmnl6HouUMLzkGfjpmHhMUKCQU
MfLT/8nlXZFnkzN9HEcpBQGyPsB1IP2UPnAzGqxr5Vjaty6OoHLi8PEKXWF5vv1duGs6xeV9HIaR
Fz1NbazELZwqnZgmoXTV8IzuJK+g3G/nmXnxh6cx/5yPDppT9ifMluwCqEcYzYlF9aOA5qMcUESL
Tqx7+5jMeEYZp3af34QjGOPZedHqTQt2gSmrvHoF0aPLkc7DEt4Ez/dx/SEE8+3s84mS605Rm6Fo
trYePij6PtlqPd8ysaI5FR/nGOwBRXAnSelUavE5+fW9P9HH7xbyd8OAwSIjaNM15pZGPSKGmOBS
9Vy6PYspmLzv+zM0DW8OaLJb9LxPAjWdRn3p49zgfz4OVByRZ1XuDq2zplUQ+fjXwBp8mslfkqM8
1aJGdrTCbY6VtVyaEaODRIv8WRvD2YMutJoIZK4ZPOfsbF2j++Mtp3+9bmXz7xf1ajOZZZt1UKrJ
rPmPHjK0UjFjhB0tGKOPc1oQGI8vKd0tC+ezi9D1SUD3kCAzhXZQazHpl8sPUuARcfu2/tJKonoM
nmdEFPQxyP+732Tgd5U84mCe8xSOVBshknVDhRyve0Io3dkNDkxB7Fywv9yI9S6mzgqMMXCtKeEd
h7E9HptFXpD6nfwZdhNe7CTMI2yhrvJg0COPb2GV1/qmlhk7xDI362AgL50jn0fLgEgshrL3i3WS
M2tc1ykw+ks/WZUe/ToMOplNyAnSEksMoR0VtpQB0d36ZS93800ys9J8UdbEDBuRSuntJxbsO0F/
C3+sApOrFq5tMG//IDd6/q9xBp8hHqocL6ZZS/Us7rdhVhxvTJw6ValiqCXE0AtZd3YgCJxb4rKa
S9nF+90D+e3fbOl2GxnQHLQRa7l2kZxVyauvmzn6c3WS9EusPxXEVHOARFBR3A1dBv0ZrwX0hnUj
3swat63hbMRHAKQRjnqGAS9DN68aiIJTv8RBw3cDfpthPZRgrMAz/jAslwdIoUIPgjlV8cLI1aZW
A9nmR+AtkUqwmwQQRmbDfxaURSfXhZsyFEV/JaSsABNYQAoll75HnQbyHQlnHqOuQcRVF0nhGWdX
qIJtsCMBTVRa8PHH9j+NLJWuwZLj6wPVSvNzAudfCIFVFJswD7b9WIEXZHD+PJIEwy1/bUPjG6iZ
KtjMhiDK0HrbMHzglhkGVzQPEr4g3gTXhg2vAuTR96PqmILTMXlzHHk60XJdmjWwzkTp+u1Krhx1
rkfdS8UZD/8aWVy2bru2nxCddabU43vAfNtHS948Prw4QbqG2WgZ3buhq5BFUv26Ffg3AU4F0X8u
AL12y8W0AcEDUBjjm/cpt2Zr2o4NLjn92uCvQshQRlfF9QCltwcKM3nqjy1XFZ1qqekYmBbT1A3H
SlvVflQPkqLihYFZOShDGXdbqSqstQzPaQk81/PT78rY+Y36xnpzwrha2RlUlroUrLDhPi9OQoPr
JFDhejhgP0mdwHCZDLjkA0sHQ3HECidhFdxmOk9fSm8UpmhSbiJB40ujPMv8PYu8kMahWSlXJOvW
uIiSAbbsh1XFZSm6+TUuJtWS5mWb+w0YOSRgE7sRPhQaUecs4BNTAl/WAM2F37x33pbC+Oz6Typ2
TeQlmWagqhgZnhysAJT7JzmYTfXE3vlCo08kw/T6yiMDIXig4TWGx3xNX/G9kXOk8G8roJ8vnQPn
azk50ihaQoO2Bw3iBDMZ6B51KG/be65vu23jh16Lzt3vezWlv6ttCIN/eFqWnbDqeHIRDvELLqlR
6rmdA3uLQyMhHLVKEydqFwNhrHRLZF0O1U/qi4QtLXZK9IBG1wWDC/Nu9V6kwTXinwKn3020eBEZ
sdkTiDTkI2v42bZITq7BGkirC+PFjJ/UNAA7UnY8TmmnHk40m8E9+mhCYTW6DUTvJIj48fjkO4rE
3hR9fDgCNG1fa3eihgPD5Tqf+IIx2u2vvco4FdKG9Eb5007wHqKvlVhbDc6/hZs3kyaNATEZy76j
nefxXDkL2GcTHn5oIR3S969PghL2CwOm+O1o8mSRbilQ6teTaCaSw/etl4DqE86+qd5y0qP0V3Eb
txa62n0/yfS5kYQUFuuWzw62eBZ7W180n8d9ukHlmHymcds1BLVulHx3TJNwmkhpCSRZBh1QPuCG
yRyWEhTM7yL5bEh0yMme2gvK1/3PWy1Uy9AWLeqlt1ohrXkFhhII0vKCh2b52l9MH0Chv9I7+6dP
zTfCk2flOIz+uMHzpXF1/qk5vSpUV5LcuA2s6oGhciMAopNiO0GCr44bxVZbcDlpo2Ry18gDmRq0
rloXvEEp+e+dJihlwF6Fn2ivI7Bzb+CO3SII5UjuWvN4sbNHWxal+QkO7Dk6sgiygiUvq4IvkoR0
dn30Mc8xGtC3Yg3YXs2EQENGiDjT84wMZFyki7/15U2mZPmEwhlOb52TNpon/GJANYgez+TZhsCX
Ady5J02Q/OfvzwOUqg9283YW8oB3HrFKL/snF85iHunY15hxMX1fv4gVGgIpOWwc+PY7awsmuMF+
UwButK6Bn2exvn2vfZLE8Ss2K1LvvI2FDOsWuP5SO8U4+ZnH2UeQQQTQR0iSryI0tiVoPmph1+RC
+Urc5Nm/vpkJifD4iLxQ8sWGeD4YXzCdQEdCGJji88iBW0j0WMr3xIEcYX3h2LexifW+dHueCruV
XHka+/G5O5K486yFjkKTRY5olpT6KkjqWpZ+nIODKdRyidEq6H4WR252QM54zVQfU5JsfzsZjaN2
0eiH35DPaIjwD0crzpgKhJR2SiJRwusMiMCiZhnDoBJReVXDEPX4ppHdBUIgpFEr23OTBdl7frto
Iw3QCtMBm4QzZ7b1jqAzKowuLLF6+Cv+sw7d1PIv9oC1v2+AKTvfxH62KZevgVBIBqYbWgxuMfk8
9GohTibZzD3s6usHfZiVQ7GqFRC0i9kdtUlSiKaGoPieF396NxzkXZq26C9+aSMMI3z82tf4QOBk
inzdFyKTCVfQZ6Zx6CTqtZK9128kXIWv2GYBL1k5qMYLnqDVYj1lTcdFOS1iLzup2B5je6vksXiM
xxUALYOactoblvtnRRi9GTSDHjcoyTHrioQHcjWPPuCLHvbnGxNh+yIQ0Rh6LVcF4477Z+GpWhln
5lfueqVdtwCxDl0/0KuXjRXAwlYdjhBvxIKU248HoiUcCpe1ctl7Xyxn8Lr+XQ0QSyENCJNs24PT
bzvkv7vjP3bZ+dY39/AgxDxrj1CJnp+mQHyOjXBXbfnko0Nb6+SUKjFw7Jhlr5QIKo9V2QXX0M1x
ep+lcSqOCg+HTt6SiFJ28wr2yar5Eyhh3K82je9cn5AJZsPqpE6NcVKnPeK5uvqO+mTsX87MyNdk
Bt4U/W3TYy9bXT7JL7yQChQWSsKR12vqyvWqNniuvEKNfmN/yrprxZyhuRGh0J848bt/FvWwpcn8
/2+sr53t+nKZFmPlHxK4Su+dOV2JmYSFnApI5DDveRmcwSm07T06KaLBOm6ArEKpeP9sOQpVEiY+
ep5SqiGdrEbtl+Nzk/pvPrsRbbzlj/EVBaeLoudCFgv3i+zXS11iS+sNom9mcYiL4kqeDl9xVp8j
BC3fIxOFbpc1s7uXAEMWn4QZGmz80DKjICo9wst56PWDgKH4/F4QZFrEWw3Ew9mFxApyweryD7cX
uoeYMhdhTd4Ldq2zuT1/muenIvdPV+n9smJjeHPrmLicQXA4nkm7jPGUuwdWNbK4Tz/F/g+AsFou
r3ChzCd0NMZJoyEOJsJmMVpZ0xgLuGs6XB3BCi+vlzqWCDI79V5m8aZKcslUaNufm2jMJ0NE2Xzz
cf9tDbRZyqu9ywt+R3iYLoJklEgSeNXQ5S9MXj0KK/mS++ShftkUhMAqzDd4KBsfhpYoq/e+zCqV
kk0NlxarDT5+V1zC4RU/0BFhasNW6rGmlESssJCNOXopZXXJIgdO/BBwxvOlBvIOobBxTYrL3ZeH
uG5UP2RiQfy5TSXbnv/CH5vB1waZQkZmCs8/poGfrYdC0BFDbK5tjF6zNQQedwca2I5IYIRxmQf5
rwY2kkQ1nBAueu7ZKknw60PNEA2eryyaVuWmkIJVrjRRSH/2N2IBGiLg19Oxzw0U+IySCU3yYAYb
i4pkilDGfpHUdULA1vuRz69Lp1Bo/4r5TspAsz2pNZkFYVYIfrv9v4axg2pyqtsgHfz/mwX0kcwi
tIVy+MLpqL3FqxKisx4EIjYfL0FJqzlq6yN3JBl7MCb3MINTbrkM0ck9D8g1tJw39UIZydo/R2rv
Jy4Gu+Ts+TiQXYljSDT6aTQYoUNA5kdfxJJIOcyGU7pNU8wkQkUrF9FRefmgJbL5wga3KEvWMFOd
PBFgSZM+N4Ifrx9OSOpXYmK1G5hXfrRK4TY2avv9cLCOFuHQMijrUJOL9/9PM+7uKPWSkqwdKCQD
iKxaihvNia5Obd4BVLkfdKLhGzutatK/TQR4bsLmNjF3Kew/QYlOWZdb8aWLGY5oe9cPRP59t9NJ
Dp5iqaZRTHZGLZbdvMT7OLYz7qh7wx8A1i+QW25W18fEGeaL1A79xISC5/1JRzv2i34FexwQjyVQ
y7pT6J9AUUh2+dZXp9nj0GbvTfQUA/EWb+eXHW7/nZkzOglYjpOqpkLrPIXDNujl6nNLGJCOfvpy
PV5chfHpJDb+W5h7fanKAZz7TKRJ/YZL9YHPrxcXiSTUBnOSygaIyQ+QaorVac0wFKVF0EMhIxbG
d9VlFnkBXtzRyglvPa3orN6CiqS2Y5tZQNNKSLHLxpNk5waOXC3o7htwG2KeWnZkv40TtC9+5e14
itQTfg/fMu4z2cSk/a/2gUWVSM59rwlpM4FJINTOXkMqKExW2yb6pMF39WrJ+40nHp7oVe6hWGIs
zrc7m6AsSIM9zziGwcWfEjInzT9bNwMwp4KSqZIJJRj69eAKjrSS+X9n95nE5FyRZAUrbPyNJt1F
0Yvb4rzO6f1MdyH1ayQ6dPtdgBN/9V2E47ZrYy6ZvKZWHI5zcnQlIJL1346qhY6TnL/Oo+oFbF8B
DR41klmqKv0sQwRB4ZV6pEgnP/z5AcX4o3PZGEGW7v1UW05BdM1Sw4xQUToVqdC210SAh6Vqk3Kz
Y7VlVVrtywO3v4DNJLgDE9SOIHNx/FjuA+ysjiey2mzzGB88yuYcrKTbvVDYsk31I/qdiBTpsp+P
7+Epa+tx04ps1B8YmwwyIYA5yJqTnqjEatQBa+PDT6BRlfwbi4WIfzAibIxfLeO0lMAdJ2SfW9SY
1U+6W3Qp2w62/HPM+HWsS3IvkfC9cfI9vvCkonJnF9M8DTioCnTkUx055KNlQubWA7daWfvToGk/
LEElio3wF0gyS9qp3YJB0nQ+EKXac2dBXjfoYKJnC80RUVYcbcgQzZdULn26UWdEMauvgOoV9DKw
vzSQnDz2mC3QGDK98UkstMgyLBkkLP+cQorZz/ezbTMQ3U17igpsrRTay69Jk6Lp1A9LaOvBQc4w
Gz+n5SxWlhjHGM7T1Az+C7oC15vFNE5vsJ37VvEeiwf2thntFhlNHz3+RaeUC/nDq5cs06MFqtBj
XWzcfufe52pSroq1I2EVIHpRTu1tOcA0uim/DrC+FDW5/bbTYuSV2zhUaEfJDP0SG8EU3+rBZ+MM
ZdubbuMGOV9obILxEqo43e0UyqN8wlFmZbFPK1ErDK6rDMP6/DdTDdviIxY+ZjEoZ1qwL11f8G5O
tIlNYllcxJnQJzs0voXaS8LHfVCdtxiE0OY95mXisolkcZBzVJhrIQzOYtgnU6NUTSUDQHrHbHKn
ps/UUsQo+3tnEdZKHEf2mAnSe6NcAq0jrWA5z2Cf95Zb/2Jl9OKAInBTPyRbYHyhBVNPXOEq/3nX
j0z5ss5bINbGv/1wzxm4RYuHxgSTFaRSSFS763HI8Csr0Zk+nad5L1tZE2OO7oGzirZaEWyxjH7I
Jr8dYCaJEKD3x7TwBk65hZFgGYkD4Db6y1c7lIEbPlfjUBDWzTkRHJj2HttTpGyC5wwy87wjTZ70
OCJcwvCLkn/gp4aSkwOiNnj1yjFaV/qfGlfKQ935HD9sL85x9merNTFsVY6iJvJLi6sU0OK2xoB3
A42+cfuOsyhaeclq6aZYDkio1NdmI4MCz2BaSYQ1yJeHcVpfn7igeVLauPOgiFk7q3UsWxqlMuHR
3n2izLZwpQcqYbNAeygyctb/nGxPiAURw4S+TNJfmELnwBzPJ6Mx6RKYcAKa+yMfc05YI1oPjwD8
JYGuj5+0ryfjb5/0U5BwHqTvJ5fTJkEktNnbfSNp3gWycrOJ4P745vEbfm7wPowJLSEOvdNHjqW1
vDwaHc2om6BsGkwvkbg4IAQ4Mb6TNfSNLExZdaaAxBhEvUka09FQaE1P53GUqAixwa76tWnQsoxF
2TeKNPUUg8GukAh4xokThCA5VLqyXY+m3Ohhm4a2xVLI6i3Y9zjyJhwj1uadInu5725DccZhcnVF
eL3zPaSNK2fT1xFhSrSpNpDCCEauLSR1t2osL6B0YJOHnYMXBkxK88jmL9sRj9QBR7kJGdtxRvCC
lotl6bN43J26aK1jml4fqqM7CV9Ipqn1vWuw1mTx6d9+i5TYHi8QAJx5o8Uw1KXlDixbCQPCB9EG
vYICZAl8QxP+maWb6NsIVtkDOmvH66Vdd1sJx94yc8XcQRu9Or4NQDU7HJ46in82fwoY4NGWpgPH
L90p9tVqyGNWQOBjuuvwME0ug/n4uM8v947958zhoyOACdUtLn/CUKnKJFrJBxlSSebYjCaFegXi
8eg9kBvUJZAbZDjpu9U3oJxyQrkB1mXd2/6Ol9fXWTLenyptrTgSWw319jCu8VL/beOGHIxW56Ls
VXAhHSpFcSIpEVPAKM+Uv8oqfUGCuk82HN1zsCXp+TBMs5UC8dO6Q3Z3NFUVPzhwtzf6Z5m2TdaU
ReaDsJKvRfT1W4GfsOGK+aXSbYGiRbfJJ5G/axbPUZ0iMx7qESWMiU99LoZdyzQSNhbHfq9gnoGb
g+1m9vTxlT5GQtsScoU7XJ01b7vkaMacGxobYnVjhCAgqjYeRbJYmjyh8N3DeQ8trDbASkPS+9RU
zpqlD1VI8nDdK48sDolKokQaN5m0vvL87PvzBsGMZAYEioCbaK7JPC1YJADP4Ir8O00Dbc79eZB1
oc7nIBCrKNHG6M0MxbznmdjoL7qDLGozvV3tzrAuoMvmZUdcX+GBK2iZbeipo4F+PDe6t/D7VTwB
lHUnSJFue/E4LyVVzBp4GyNXvwr3cl365bO/Rz1rRphYWdXfjC/UlpjVRgwAkz+9HUiv3s3Ot9Ah
A7aRI77dVg749LwHKCrWQcZi2j0U4WY7v17QtgesFVu1jc5bIv3ENBH/noFaLtwedPGa0nPwmr3d
Se+kSfpZuBM+yT6MfDC+Yzp5fhvek+7X9a+/ryw7ZNnHEyz3eNAArdf//y89RhpFDcc5T74T3kkf
Mn99GyCC9ji38DsN9nv/Kw5GbnuABcUBXy61QOQNToknmEKwyWT5WEqJVyIcWCXeq9MKTiQ61TR5
smDu/v07LYesO4OehinsHh+bqwD+YSvyyfmD3gZd8n8FTEbMyBmj11WvwbuL1ROu5ve4TRWeYPhH
oJfsiUu3QBpryVb1/YrmDY2VccpXNxHCuTXYpmH14RQOwdfCoiyAJOz2A8b3SO5x15Lu3+Gk3Qmp
L+4DjIwt6EV0fx0i9N06C6Yu+lUlKLbl3/p63L5AxE9pA5gLQ7iKHPSK6Um4zfInJPpTqb6vCFn3
WSOUYi449fec/FS4tL8Tz2GXEzhK7X8TB7bw1TyqJZg014vobiI5W7A0gZAMccjZdIJAPZm3ZvWM
1WPXZe5sRyjz09/GeMyrSprWzqs2EAHDHRNsJy/smDXFDney98c4iMPfw6cPII+EGwnR99nSmlOF
nmSVV9NFG/TJ4nUSSxLeZZJ0l0Cl5rexEonX03QSGir8PaDe+5w6dW6d1DCDmdV9aLHxrCUJTJoN
eLpMvasS8cKpv6Uw9sVgmHAzikm6oIly3bvEfppMvszZkQsjQylrFSgQXBViNl6KvZsnf2bpbUTo
ooWwgCU0vrWr56j5Yv1GJzsPq3PZkO6icdZOotSLfLNqZIu9kAhvSjHNchpNeM6DlGhooSfYekQA
LxY4EASsa/wBmZ5aDh2iNniY/A73j+utQDLSf38Vl37UrhwFyZpQepg9Q+It8MyKdqdNckke7nBU
uXsRkl5aIUm2UFM6Fvw2FhC2gnBG4+nlhhCVmboJYnXyXNsjvcJbmusaDm+KPCBR22m2JTDhD9Ej
Y0uhT3FWZe8sJHXycsNjmubfrvCKiI00Hak5R6MpdtzbXZcqOqgLd/xfSUs7nP6wE7Y++e4v/g2O
qNjpLz/Egtg0GOtbeqP57ZhI9lPWIbcQw7yc99Vh9GVGlFz+oosiTo7wHAyqy83RHDMKyMTy8dZo
fofXOkiVcZqUWUIfK5pXNWAh1XAhDdDLnW7qzKt3g5zvtEM99bv14tSa8DsJU/sqFyWwCWivo88N
UQ6qK3HIGHayh1b80fr9JSU/PWENtiSRlGVf+sWpWt2Ds1GpFs7DKMGsU0RCuxdCr22yctrAlQ4H
RndltsPUClFgM1icRkHS2BO0cTTz8KVjTz2H10xJZrZOk8NchSLT8grosOEe2F/B98equ9pfMgi+
25Ff+vYeSVREvkgiIR6mYdWhv80+j3H4A0aATT3IAghQVmjiuYAm6Z4Z0vuzxlNhj4rAynd5nccL
Iz/mWGmWvTycMU1t14TLvkJZyYD8KMdOc+d/EYErU0gwXzt0gk2mKXQ4LFwI/w5P/BPeESyqLi2J
vGZx/aXQZm1xDSSj23TcBo93jie3F6xSvj2+y+GJMMKZ9215cAurUAcKZR47dNrvKdVTNo2D7aO1
QhR87YUquX8pVzH37tjt6vptuyDdvNG3aV3sOX8cjhNSmoTPLhqS9WNsjsLCHJy8ftbj20VFjtxa
6R/e+nlD6S27Th0dhHTpIMri9eSs56qkA+mgjl24DhYdW2hHUwhTsPZr9ZKngqW1D+XgwBW4oGtT
S3JTY6ZuBjUK7LaJ8q+yStDD58VrKo2LFlNZhvIcsxWa2iAC8uArTCSpIOqOE93tM+1aD32BXY+w
DuN/ppW56106h76LqN1e1ITg9auZBpyh8wejPTXomlzbFD+NkpX/iJjKSBK0eEXptyAaqZZHuyXN
fRyqphemy4JeoBf1V/BP5SVHDda/WGc9nkN8ahmyNe5L0Gi6UmbWuVqTksQ4RU0IjU0Ehq/amahP
lxcIJuC0TPxFpoc4dkoHMVi9XWh7d0DBEJXGJSHhVa8y/lRjjrL1gcQDYYt0xxabKI6x/m2ZFdlh
scLJpg77ynXduGJILdauRwpR6hN0iD9bzz0cD/ViOhe48vCC2FwRUv2vqL9Ar3zDkYO77ansFscW
2C7D49h2JZ0Av7b/lPQEe+izR5zovLfYcau3cy5Sn36Jg0r28+Oc/wdpiqgIw/UQoZhj4w2/T8B1
SSzqpuYlT3q6jqA1+nyVPpoUuAEfcDiAeZNz8b+yOXBM9SCM6/nKxvIX6xZwaN6/sdrAREhUeK+x
mhj09x8Mv9LZ5YuvRX8OxXN6KNSw3qzMUDhYP7vJ/tvDFc8e3ySONK653NcNkIPNKhN8uhGJ94B6
eBG6mUEHFwyw96a/brro6YsrXbWi7gAZ6xEmQ+6UopkmiUhWlZnavZUPkO47bEGTkugq7dp0d6zt
7SYTOP9g8Y8S4CkAN6wO8Uk1EwGVMFNOuGWle7jHWQHXVkskrrDq+qOe/0xaPsso2halHtA5WZG/
gXqhXdO1v0/WRYvnJx3BsYsuQICSYIh6l8X2XLWmecluMkM/8SRtnLi6wJRY3AHtRGJBYFnjqX1W
2zaSgjc8OJ4bRbu0OKetodOSplDt5q3CdJZCD+C1JT6T/GdIMSsra/MWfOguPGY9rnpvqjkhyy81
Jt9+2m6uERB+ayxPncPKqiNxV/GVF2LVt5eXBb8Hf3rtrt4WqsyW2Oz6vy5KF1lbTrvYZs/SGiiD
rRe3AEkBulk4ZWy6DHiUOLO1URTimW8CGrq4Ztvk3QYq5+lv9Kh4OT504XGojSHW328Y6uvC5Keh
fLCwHUST0mbCkI1W915bkuK6Gl3YhJYNnGDdwv7H6xVzDc8UNlAOi0+quOl0POiLASo7Tskuhb48
yWNYdAVyEJDUCqBAiDUUPg3Dwrr5Ui8zGkplJxbcA/PRBc1GxiVZq1cXeTCyPqgCFy6SaEx0odxc
Aqtk5q/lNKgU5inVrl1ElzrMtUXqo4WSbJwJDOzH56aDQxC9hvt7wrr7tJ82rI5ZCMQj3zhT+enI
998aJ0SDC34WDc8I/3scVokw+U9cpT5es3QN0uuZ/BnRYkjrylzahQq3duDBShrWrOdKzNJQK3b0
XcyT4tnWh8IfQXcvoMSWo3LLyFZn+VwTQdw9o/tZgjyGGg9cVF8+ik4hwN6YBbTS+qDQTjs4oJA1
bgISZcoc21F8TOkEpKeuSrIlNtZGql7FrHHuRJJ5j9wGfcO9wEZnQeJp51V/Wn/Ba9ol3cVIJ9TB
QUagOwtkvLCy0xmhc1r230owN5Ux/n6NMmAra9c4sUXjirtNAI60eIViM4gk4cOeS69FITeUVcay
4Y68fuCe/7BiLf5G5nZzN0QiKfc2AMjL/rv2vsVCpQMsnqzGZJtxr079G3+khdJX+buSj/YD56Kh
787Sb2wq59c7pJ5gSyUUGdEnPQEeTnd9XmEsOFAO/0OGwDl1nMSvFYOmUtL/wdb99lNStX5/cutp
+rfZw5JfturOtL9qPrPrR4gCB/OzNoDLTfqUiRha/lVM1oS/WluCLTOjDz9Y91EVkaH28R5Tdf8x
4Qn7FRbPgAmbk+1alnF2byPw9Z077FeQI/K7iNGuIqOiqNgD+mtF2hGQv8IO8YS2OiaRItcHnY+t
pcoWBQ3tbLAmKgTMOf1a7/OCIl+8G4yQpPnrVdlbIuDMUmQg0yc5oS2laQ+ob9zHH10nPgsmJ1E0
eyRPeBjqM+wFQLq5rXB7G8I3FyTh2JoPLubFeNzZxibmq1+YEtcyWoXOTzFzIcmhkGOxDTrrX9ce
tHOZFgjnw1x+66/IhQ0dBAqaGS6+m2KpZqMJst3kPUtzc1/NkXg4r+g+Ph2/eGcFnYwLNJ481R99
Rc/63GsBoq2UKDAFe93S4X+HDwWxrsFFBhYMzZZohiICkqP2oW+M/amkqBKKn8dP9COEJeuv4V+x
oKtxciCQt4gIG6ds5cQZGs4bH2j+T5GYdqN44uUfgF2GKQwsgR4A2cbl1D7uX9qtLfB82Dx9yxpN
EYNX5WbjGJyjEWsNoj8v8FhEQQGCAbx9ctY+33WUmH0QGVI+U6biMQudNakzaBNxcY+nXl1RmPz/
eVosAd97L14PAcjp+3onMBl4TRh4367uep1k386zh/0XTa6dWB/bb5ES5aINrF9o7LvlyvRerBCE
rqN1ftjYbTn6UDiCHZRt/9wxVgg1Pbe3jNWr/loLDnSflrtIdQQzx5yZsQM3MvF+B+boNrUPKRQC
UoBOXXqG1TdyiKtzKx3nHG9Nmn1QswLlgCnwmU5EneS3k2ds5ZWbqyE4nESSFNuLpw9rDXo/hvT0
XTuKBpybIkUBCiLX30dgWLpsI69VFCUPDJB28/egxKaN6qx+h8JFM36RNPGHcp3guSMBPHGJd0I3
97Oo4BXUZUEsLoVTZ2LxPiptshbAStTq/j/LsBrAB26/2AkwMvZhVTYuJ+P7rTs69/Bx1c5AWbQd
ms3GE72h+OFIKGiingDGZqRBDTjvIBspWwb3HaklcNzI6XkwxccYEv4MUBpByGVhUMxMXG4ODha1
zxBf0Q3QYrL5uRXc3hOnXtpVUgd1e04zlJoCk2ncSUF5n2iC9ftrWW41MfdWokxXPYkKW/1kV3yl
DbF/t2vzWp3wm3A9q01K0xuAuY9CL4dZVCHkeDEQRZnsseblUuTYO3arOA3hPEMKw8Y03/KM9f2O
bUjn586t/vwPncb5GR1GMv73kVCmLR/wHl2npFyblk/iBkgHa4OyIoS8wnXM4Rm/7xSNbZ5Ffw85
RD6IxcqVeAEYm3RWYF4PmfLh1rCs1IjQkW16oSqWg82DRoKJ6ezmiLKPHVT7Ws36jDxkADjPpxLI
xH3dl/oikCIiTNmFUaAbAxzmwh5lmxsozR/3ieZmLDTFwM+Z8uKdOj7yPMtn1M7BkLThZjm+Efqa
lHinP/v/jhCI22HGc2zGBpEOlxcULC6wpHcGlBSB0EhIMwhelwxxgWOfepH1zynqYbwt99wIkrmv
sGRR/0/Mn4FS5CBxzokn1QdwCxtQK6lswohtdoeP1/lO/zvJy32TayCGPrFoUlvBPEvp5NA87SQb
Q3jeLSy96H7JZKwmH1SaI/9HC2NyIUREUUQohndx7xohpKqQBZa7epnawVymt1VKS2K53CyK93Fj
V9rNHCUDbcbMup4nBk9hMBQ+jrBae8mHI9mUIiqhTkYMErwvaJXV3TfFSdYgIyQOSIYkxYkAirvC
5FpzfnhC76nKFUes1k6mzmHzuP6e8nbXb6xL+lc/wlUZScWFfGipaEc8BAdZEbXfNKwg4YyvpPdU
wr1K3H+8lNv2MEDS/hLMWLQ3Zprn/3XEjt+vEc4fmTIxg2ZfeqkQNgm8vVNLNiTQ9PsUkNfslVIy
rvn1yJJ7uTOrfJq85OSfgkTDAWb4d6nyCBPvVaT+Q2TtZHUNagJ/TB0cl/FapnIbvudBpEWD0z59
9HKYsogtLY8bwisulSqsUtBh3niMF4vS2xEfHN5htN2TKd2wYzFF8z+eoMl2eqS4Zit34a5wCion
J7KyCdmZs5iXXuKEmlrtgEFIHYrRlAErYPQ6Fag2bIXXTM7ZbfyG4tFFntiYkODuRlOGItRe7FxK
J13oCjXnt13iN3r1x7UNtezNX9nsfDNK/0/Pc7l9rYmZl+823p24orywb/vJPHEPWkyxVuxFXGIw
dUTV01+xkxj11tHUiqzZyGBTWckAKBPMSbEee46JQwOrFCYw1xPqSLahN3Ulf2m/e+djAUk3hANC
CyKgxNAnCdRHevO5dkEvG/p/2W/g3tpyLJGoMwYhE8JF2JcZHkCItILZ6GOVxUiDDJbaE1VEvB5y
owGr+h+AlG013WcaHVxss6l6bxtbz4HD8favRSVddbZkHYHlZuCah55jA88iSUv34XOTRRl6y/95
uqKJMbXv/0ZDds2I0c2CZDlQexXT2T5glHsvEl2GgQGAnHQrwViXyhQjB1EJCmyyyf0E9yePeJrY
iPDLq9GBQzNNrFSo+PL1IqzJTH6oOQQDClwbPzb0xtlYbGjZ6Jt92KyyTrq7yWtucbCb4viJYISZ
89pH/g1nN8yCOOkBhXHIUuzUlKKnU0wbUjdnPXxOecD0tr6pv3jLgSXoDgfv2ONLlt4EIBlZQTJL
jhGsxnEoiYHm+91/TlutYnjKbaafuXHeGDsZ50w4xJfFBjO8sbQDVVvqttN/SWdvrg4Y68K4HHyR
8ajrRPb5kq1jTg5mhy/tYDnqW9yfdK9u/on4QfoJy5UHv22PjvKUQtE6f+UxR6/cum4TINkGdHXG
KokOgK6c6e6d4GZh3FAKNCkyoyN4LDKMO8eqh2f/lg7+F7Jivyh4t6OULbwNESAjoCGOr11kyNxE
7KGL4DmUilw4yRufw/n6vr/qW3FnVrolWv/L8bCkkTKnUJsuJdH5RjbeYC1rmaQUjH/7BBOAwX4L
b6HZMOOyBdP0Y4P0hepOdZtoGtilnvIpqrASx9bmIKAjvhZrzdlsAIvUry0Z4DlcRDd4ozOtNE5i
1mu+jnwRrT9spbsSwMtO6GuIMXlNDBZrILn2//I2yRcsopwYIuKLJEWxDW5OjBbo2N7RO2pm2HlT
2MHEuVbujAoFc//as3hqkVciATpCzg8sEq+Rmvvctsh8iGV3tX2iU0Gaag8WyQZX+OZf8iy9gvl0
Nc22TmTDbtrQ8XryGpArVOmbz6mKr4p/o5E2C+ze6M+UHhLeBK8KDl6WD83dGKo+4vfyTMJxObv/
Od/C1K9pzZmCJFaqIUqC2ciwAYAydx3+Hx4DvXsXy79bpfEwdMJTzyVkJdgKkLc9edtEhkB0J7Z/
0PtrAcmfhJh2oEeCxS9gZJz2Dwxb2ByTw98FCfeh/50HUAc0WDUOm8c+OGjmJ0+y2ibVpqv9fIG7
3WGpLKaI1s8GmptPSrqJLYWIADk2exj8Ib4LWT1BbF/nKlgllQkX6t5LYjduoKdGJ0e7e0XblErL
SvzggESuQWjDXswOuL+4fPoIHnn6zaDPEpzE2DsosEBX8equsYAd7JoT5H3rRswz6K0P6Mn4SYC3
RX9uAEWK2noLCtYdB/wbRVUqLp3ZUJog6PIuxTN5oXuvwXi1sQMukeJFp7/SsmZk+REWqsw3+21B
RCMymT6Ipn84ouX0HN2i8pUlf7Ymm1VGA5XSAFw4fHr0ahNpmYJf+RTGEOhYDQKYj2FjQgDg+4pW
NrwnKQKHxT9Un0XntRbFSWnqh89XZmMZnXIQ+g2YD0fgoITNrlgoB3m0gmHx1k8OpAD6UqJiFZ75
GBc0/K0yYelPqV8/mgIvOguld5x995GD6ZO8uC8DkEOENh6j0uQvoNr7rG1gSKcES/T8GF8crDRY
e+Cb0aHX4eOyPDEb7qwkLLt6lwdWveaw1crtjR85eGWI0EpzR6XK4XT3r7RherQpNcYKnJACaVvv
7cNC3eXTOgQfqTQMU4i6tMHkW2K4i8/qbyws4lWVOGYCMy0yy1FzdIDCzOwFcTAex+vnPjlDEzYS
HQRE3Qli3dXYbMOaLDcSciPQDpFGgd8RnCN5XnydThBKTRtuZVzRr++eScis7ETzXmIUzxiwlKY8
foq/2aXccNhkyfBS+iarCiAIqqLuB7NWnAfW2xgiHxd+tnhXns1VUSTMujWS9yy6mf7y5Dktnu3j
kmYuH8Doyr0QImCQNHtgWN6AiafCNcWrN9FqzZubAA7J876OGhIZ3B7h3s4ru/gAchipowgas8sX
l5aolyZWqpGqRpmnLioYoqAxqzlN8HjNoUr4ROpZZHu1ujzASKx6bP/IRPEDGmj+g1iMbwUz4a5y
hxdnYlQF5eUsrJ7qSJTVeEM23oISBfzDUGTScOPcBE1gGMFowTaYND/rcL2IMW3DFy3whlUjYTzx
9LYeE5YSUmA/ZgpPnd2uCPsokaLYMAcV8dCVvmdmOXo6oQYvpz6wB7jiJ8acEnYMpnX8aWRVPZ5p
4jpuVts1lihzLsK/DSuSyTx0ymp2oBzvuEouZB2IR4GcwBoyNb4J6YSDrWawb/e12Qjr4rg7TWRp
dshXomc3q1LvM/E1G7sP9nJEJplpXjc7C/5q1v04x3Rt3NXDjUzKbaLav8B1z+A57R9i9MVAw0n5
48tMS6FSxmcrk5korDmAJHFvaLOQ5m9NxLNjHYMeKuhci6a3SmekSoEHmJTivNYamS0XTIDxo/pB
UZdH0hvPne4EYL7ag0b6OK8JzprWyPadwJnr/yxJSlZlmbJ24+miyNZT1z3/bekKitOGs1bLMSfA
8hlo3DdIXO5u+F/KoDkugPEI+UR+/hBzmA97BvOV22eqhDbq4aMngfAAID1M7x93oLL/SBa8Oz1t
UFlMJRAqYTQIg5PrEzB5A+nx5Diz3JI8XO9H9clixtAFzRVEda7dg6hn9MxnzJLCO1mdBKQJLNnV
PmLBC8grlgdIiBfmTEhzudxWiaATcCg2nFSruUW3kXOKH5SJmN5d80cguMoRkFAjfHs3v/GyX1wJ
5HGF9CZUe6phqgevX6iReyFIqxlrTbPhCC3mtXjvIjFmqJjAGyxQu8X9zPuCtXJxdOa6B1QLV7W6
c7CLRItXbocRSQS1M2/shqoPrtg5XZSdTUC+QEU/xUMljjZV8kq95lzgeiMWIBXeQLeQvmneUDX9
60sClxOKiIUyE6to8ZLggOGUkvJSGFFB9vVdKyO74A/fkSLT4GvyIKPllev0iEEcb6MuTX9/4OTm
oa8G2f0ox07fKufxtelegTv7EPb9l6WbyhW17Tfu3VSMxA7qfLcqv5T0rbv6jZurUcl5IRbUPXBI
sBFGLrDrIuItu3HEJoi1HI7wbQbNNJFQjDVuWlYlyX7vE2oaRhrYeE1S1Y3Teqq/MZfLFtZAbve5
PIwZRXpCRxZIWsudlJE0XvvXKPRKDNKiOidk6cuwewSqkS68FugMF/grHgsafuOJRsj3ZUMXWJZ3
Znlr4/pstQYwmHXsPmQ0u/8cCr8lembs8/OzrZKZdI899DEnf9a4PwF7jUasvE2OOE+g3e4PwP+T
3T7vQNU6z442OkFHpMvQv96VY5BT1FPCVpk07Wa8CGIJrxP9HDXkwtXs3b49LVV+Uz6Kggu4DJfb
pMH11HDCwIXMP8/rWKtGbjL1aOisrAWvG5Cye3EhkXnpWM9shYVz2IXzF1jVcjpmj4JvS1pyaSFZ
0zJe0vyZtNkwj+OG4ZuhHKLXF0yPqZJv2S1fqtT+vHts/WooFb+n8HZDIhbZv0y36aV/6QBkpP3o
UJfIgDfa2GKtCQuEQISA+pDvzgtTJoP8UYQtQ4XX8R4b/cHEvVoiP3fD/PpbFeebqVpeblRRxBlC
1GVAaxM6ggbpz65ajYomtOIgizuDdHXPN9GCGpe30i8nL5Wt3SYvHa7GRwzSkw/ls2DoNknR1IfN
bMwjOvRMnnBZULGjjxR/aY7QvN0f1jeh+oM=
`protect end_protected
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library gw1n;
use gw1n.components.all;

entity Integer_Multiplier_Top is
port(
  mul_a :  in std_logic_vector(17 downto 0);
  mul_b :  in std_logic_vector(17 downto 0);
  product :  out std_logic_vector(35 downto 0));
end Integer_Multiplier_Top;
architecture beh of Integer_Multiplier_Top is
  signal GND_0 : std_logic ;
  signal VCC_0 : std_logic ;
component \(integer_multiplier)/(Integer_Multiplier_Top)(WIDTH_A=18,WIDTH_B=18)\
port(
  GND_0: in std_logic;
  mul_a : in std_logic_vector(17 downto 0);
  mul_b : in std_logic_vector(17 downto 0);
  product : out std_logic_vector(35 downto 0));
end component;
begin
GND_s6: GND
port map (
  G => GND_0);
VCC_s0: VCC
port map (
  V => VCC_0);
GSR_0: GSR
port map (
  GSRI => VCC_0);
integer_multiplier_inst: \(integer_multiplier)/(Integer_Multiplier_Top)(WIDTH_A=18,WIDTH_B=18)\
port map(
  GND_0 => GND_0,
  mul_a(17 downto 0) => mul_a(17 downto 0),
  mul_b(17 downto 0) => mul_b(17 downto 0),
  product(35 downto 0) => product(35 downto 0));
end beh;
